��/  �Xt�`$�����My<~}�A��5@%z7�FH\�0��-�9EMx*1�s���v�G���n�2uO#)�Y>�P[!W�n)6����o�hY[�ܾʰ��)�q�3����ϺeK�^)p��Hz�{%,rU���_��^�^ۜ���l��1An"3�"�����o��LV�laD=tp8F�:9 R�ibD�鶗9�1_>Y���4$MX:T7�q��N=����w�XEE���?��&��i��(��c}��&��>aӭt��fw�5)���; ��H����Do�6	��gy]њs���Bm��.�E�e��Ļ�60��NP��ب��Wx�z��Ir$%;M�I�Z�<6b|��m��P?�0<s��w/�8J0���:��T��I�;<�l�Yy\�7Y(
�����I�u�� ,uQY��j	����6	I��4�H���[�0;�F�$�ȣ�3�+�6!�u��׬�2~���4�kWf�2��]o�*��L#��z��'ى�.E��|��s�P<,i�a]���J����~TVhӑ�l�s&������DT�ND�5q�gl	�7C��r9��x�o�cy��:���w2�&�y�`�"�����W�+�;��g\�h���Ȫ�T��9{�E�#T�y0�S�LC�ۆ���k$;���9K�Q0��� ���Ɩ�o��|4����[�K���T)0�W�����������mh ���#xh�SH�]^e�M�Ǚfmv�~��0���6� ����З�55�Ac�N�P- ���uN��1sLcb���
T�~�\�Y�4��&'�%R6hP���A5��$���N���If�3wz��?b��Q4_��)7��x����'�C�9��~�w��<��qzcA��앣#�9Ö������ń�J�OQ��Z��8����29K��"/������F�[����	6>�kg��ߞ��]HV�pG�y��	��g�G�j]�e���:�M�o��%I���T���+N2A�H?h1|�U�{�ah�V���¬�k҇�E|����r��(^�ȱ�d@"��j��S�m9��3�e��uˎ�1d��kC �)�S�	B<��fΐd��<�e��L�����t;#�z{�Z��>�w��hA��|�)�b�j>��px�)a�����a�>j&��$�Q~W�|��e1�?�nd!TO��b�Q���Y�{�)���	�e�kP�j(}�(g$n:��e
��o�O:���5�p�쏦N|&��2��G��s���ԕ�5zNV˨R�:�픖dr�,�%�{V�5R���ѩF��1�>��D�$��3dy�`�T~�b/,)5��+�%Ŀ��XO�~�#�W�}�]u'����y�C,����V�>�6t�u��� �fOt\�kRl�uZ\����ڻ���y�!t��J�s�	Ld�q��(w�|=�wX�?�2�u�*�˵��pΐ���[�� SR�UM��؆��^�s���YD�q}$��^iP���F[�0l�m��q���5o��XNq5�x�)^9(�䳎Ԥ��i�%�8dR������Yf0�?���ʞѕK�R��s i�nX�AȞQ_a{���^r*���P��E�ȍir-��ȁ?Ҭ^�#�Q��7��c�O}.Mf?��{�ts�d���5�ivC��\�l���ON���^6/�����p3@%x����/����q��!h��a�/�.�?��p%:^)����bSP����gݣ�^���J�Z�ӔNF�;�H�^���?K@1���G-U���K�l�:�ܨ*V��e�����v�ׄ>^�E����"@p�b*vaG8k���L�q[Ve2��X}��,*e�O�d��=j')^�}��U���G���8N�U�����**� nR*C0��F+u%�JS@\F=�b�gCwΩ�A�"&�f���I��5?\'Y3�ꆣ�Lyݩ���@��,�6^Κ.
dKKՒ���?�?���ӛX�k��$"ړpbu+�73�d���J�6�X��B�#��2��b
��������F��1%��Īn�R%MP��lw�|vP,
�Sw�e]�,�P�il��k����N]ۯ�E���:1�,��L�{��L#��/F�3��p��g��u=s?��r@��S�
�o�r7�u�5�B��*�1�&UYϼRd�cCZ�sJ��K�"S�>�6V3@$�[��q�������3�}j�0(�?,�M��\���+,I-M�Y7�U�H_@�������h��,d��S��w`�/�V{��7u����js��`�}x[G�g�vLA����d��l^�3<pfӚ��=ry��!aq��!f���
��g[��"�$�%ej��VN�H;��qCIM�C�ĳ�e�]���e�K�oN�z(���S�_���*�I��w����F�5��<Ҥ�V�Sj�]���3�����&����Q����a���Z?�2�i��:*���zvW��cJ�g�Y�03[P�iY�V�V1]cA~�F�c�+��9ذXF�>h����ᙱ5a�%��k�t�K��E*�(���C�M�O�cEx��L�*���&\�P���a4��m�ǯ1�*�c�("1�{[�pv&d��9['r��Rn�Wd��=f�7���� *��l1�0��~i��e�k���?��R�<kJd�G�Lh�*1c%�p��IB�?�s�er��������'(N/d^��P%����n�$�@�]�D��(n��r�j�Ÿ��b�0�G;����O�WsԐ��(�:UWL��vT��W^������-�e>C�(M羀ɔ� ����@��<�߰�����cX[��7z6�{7��C.��ntt���������y�h��>e�q>�9Pխ�Q?6�F�F�9�����YM�U�lew\D��C��B��ùв1�i�K���o"���ۍ⸲З¿:P�����}[+�b�Ͻ��jLn,�6�����_? <�ڱF['������%���H��,������}��9N�W�����RNx�AY�cɞ�?2�i�&z۟O+���MFC�$^/��J������TN�0��p�HΗ����W)���q휝,�`%���/�HwY���J���߁���BU�B��A�mY���~
��3{X���-n���0�#ލ;������g�2aUp�T�`�:ԯ6;oH�lw�r�����oa�i����3��EV
Un_A��4K[�*�Q�0ng��\�%���0#j�Ȉ�Z�9�n�8yM�����X��$��ީ̬<e�V��G�����j�#/�z���䤿j1j��-��V����<��o4q���.�Svb���LK���k���������MEh6�5ґ��q1���7:]��h��i7��c��}�;Cj�ID*�?���;Ckp�J7)���vk�߲ܡ�c޺q=|���塭�h+
��:@hͿ�r6p��b,7_��������c��� `|!@�8��$����	�u_��m���tUӢ���1��p�g����1�|�Á���DIN���Q��ԧ�U�NC���#t�6�t�8, �l��Xt��gt��&U}w<����䙍�E�p) G��b���ȸ���
lF
��{��:�h3$�o��3�8��R��\��g�rM^j�4��諃��qԨ���x��$5���c��6�e
x��DS���&��t�� �-%���G��:eKtx߷�k��֤��e� �;o=9�� �?�G�̭��Jtw9n�*�E�n����1K���E03����R/�w�(+�m�u��>q�TEƅ��w��W�n��*3t����x��Si`H����l��{T0�c��bO���r�0�H>���.@_�Oj�/����"t
I�Ւ��I�[�r������|���L�G�n;Q7�;�K�Q`�Ĥ��M
>�p�U�4�h͗�_Ls�7\j���D=S��X�W�9����I��������.��b��D2Q<���%�.��{�r�L��3@��J�q~]�T�ʿ��?�V��5�wnK�ۖ��"I$��d�տ7�/��-h-h�Cb[I8�oZ������{&�s���=u ��$R�ǿ��ٳw˷ܑw{�K��
Ie��Ʀ�g�|��#̽��đ�G[�&����i�-{/�iûPc�/(����ЌDf)��h��&z�CR��XU�0x
�dI홻0�t�>����V4�����:-r9^��W�x��7��f.9�]�<�ٷH��?@�O��6d�2��|���4u�#ʃ��snQ�k�v~�����Ⓙ7���&>�re�xk+x�/{�������{�2UI�YD��o��<>
�Rİ=��VV����G� a�JO%�f��4��[�8�k�e<'EmL ˶3����b�$���cqDTŵʔ� f���}˝b�X�~#O�#�=@�!WS�9S!I.��*1���������G��N6�ՄC͌[g���J4�\����!�}��r�)C�E���AP����y;�������1�|���4e�92�p�@���c��T��i������I>q���\ou�T��s۶�س��+�]��4�S\�dr�҉/�S@�U}�v�ɉ��>�%yw�RS�#��3#!��oUB����vCm�Ns����M˭�E�sSeGz�/��ĝi�j:�#�nӮ�Tn:B�O��1v�ܔK�c ��������VrTsV�yP���b'T�5]�*dG�帮��w@Ԩ���5B1�'�8�E��pֱ�L �8U��]����;�R��_7���i��3��:Ū�ޯ5:i����:+C���;c�^zG#J��F�!!~)�u�qV�)� ۰�]�AP�O���dF4�ڷW��|����"ٖ���"�-Q4��F@6�a[�*2�O��m(��́` f���t�i��)���P^y ̷�%����vI3�UH���j�[�L��g���<���?[�wR�Ub��V͠������}�Ҙ��L�����2�����Y9J����ǽ����O���Aҹ�_y�VB�e-v~��@1�zqF����:�� �c�Y(���(i���l�X��kә��h��7���!�Z�Qĝ��{�7q�U꿅�~��H(նD��������K@�r2���Z��m��@r�ɍ	� �A�������\�˶70BO����If�24W<ۓ��zxz���a����y�YA��+]bs��U��H)��
L?	-��t=������V�F��\^N�S9BZB�t�'}v�]C�=@���(3�G'��r��8�L����CT�؍}����v

Leߋ�=s !��r}��A;��G����G��
2~�E�*Ė�aט%E���nY�XS�y�fRo}8Rh�Ћ��l��R��E��x��}dE�w>K0���b|�V������o���4�1����L����m	�*�c���W�a�a&�8��}�ʊTI$�g�K�'(I��z U�}��%��3/!>����c�Єqg �̀~���k�����h2n�Mu��!kHVvZ�U����3�p�7�0CLߚ��B�]��뗪�ʿm��F����I<A�4��#X���|3�Q5�Q��5؃�%��"���_�1[j-��0���*>�Ϳ�S�B�r��Q|���&�L3��K5:�S�F���w녥q��$]��F�3��Vd� e��_  �A_eT�^�ѻ�;,#J����	�g�R������P��v��-��Y��i,�2���H����`�ޢ	^���]�u<��
"_���`#�<;�-��"*��6������z�O=ԑ؊�ф"]�3bi����
on��y���hM��9�Ď�?
��ff{��?��O<�`�>N��$���!�V'���x������Ⱥ�PE�%�k�<xϲG���.V^,�x��}�k���݃尾��q6���]�k�L��R!>��Έ֚�C�{6�@
�� 2g������51�h�7������<0l�7P6��\��C���g�0�-��!�H|C0]��<�O�U{A.C�V2[�/�ʪ�ᣚd��x]�2'3�qO � ��*٪��"���WxT��m������b��^�%�y梯��w[��tLGѐ���d��X����zvZ;������P�2*�����	'��ڌ=_WXY��L�*'�븐 �j�~!���6������A���XA�JkoK�&��`�kxgIWqE��ק�Ǿ9^Ji��}��D��n��!@i�*�؝�y��{��M�Ǽ���+�p�����2*��3�k�UC٢h8�d	�͘�uޔ4����f2L܆�K�#��댖x�����H�g�Kl'�;z�\e24���0�08������8�i�Џq�S6�<Q�q�BW�����&�S����w�{@�b AD�]�*7�8��>�	a�W(��Xe50V5-'�"���^�۔gv3ˡ��؇y�Ep��T��8��aI���;2�$'�:��R�F���eA��1GĄ�Q�<e'�$�wBR6v#z~��v�M4��z���%<>��ʭ�M����N#�ؗ��/�!�	�)y�¦�Kw��X�ĕ׊�mk�4�T��v֧�.L�aR{�w��ADHz�-c�}��k�{w��Ѷ������q�'���%�@��̘uNaX��4����C��
>1J*~��S�+칏9V� ��ć_A�0�g���k �>�������(�)�]2�� �:z����vѐ�K/.b��ɔ}�u��L
�,}Y��<̾1�Ly*��d���:a�-��3��t�ib2%�N��K�+>�5_�|>JG�l�3Ģ�������$.d���hE�u�V#e�HWͫ�\�yO�V)`��b�y"x�ikd���- f{u������^�T������[��\EQ�) �6�&�ury��݊6M�[�{/j�BAN�msr�+m(�>�F��N�w�~�P��8���I�̶�%��4�='^�dH��;Lzq��ZK��x�c:�'�]Âm��GL�R]�	W�5�sHvV�)�&*�3t�r��@�x8F�a��N�,��2(2اr�4�n�EFF6lU�ü���2��4#�U�����a"d�g��V���1�V��K���o�T���eet=�+���L���i�O��dv�0�����3����.�B�:������K����;	pULPlC�K��bk�9�!����k[�#�K9vO�^{T+t0{�m���ةH���M/�^칈�T�؅���+m�i�ԯ]�4TIt{����>�Z `���U�F)o�ۥ��v�F�Q���UI��jA|å�YB������N9+S� }GsZv`݇�n5,�J�q��s�C´����(]J,CB!���|�1��Ґ�(�s@0諸�W�ă�����@4�n����u� �~+�\�
���/�0K�w�qV�Ls�ҿ�n�o� f��|�Sv#���iDTt�J�}�l$�?!�z �<-Ń1�I8� SG���L	��_NP|��ǳ���� �Sm�Uܮ��A�Y�U&Vhx�I�7��l�I��Б8�c0�z�+�BD��Ѥd!^v����Brٺ�F�s�ZVK\*o�&�i"C��qne��tϷ*\g�=��3�w�������p��6U�
����<�Kk�j���-UN������@s
Ġ�s����|�N�d;+�������X���6��k87�Y�/�*� �ؼX��;�j֐���V$_5�,�gb|�)�-=>d*��/5�Rc�/�u��qp��xOf�j#@yMޓ�2?��E����3�-�0s���qTQ�J#tL��"����H�3n�6U�5I����s@4�V�u�E,��
x�^���U{_���a����-�_i�#r#;����/_3��V��������|��Ǌ�K��ZpD��7��fĊ��1��o��5�w��������Y�-+(wOl��},����:�z>ȡ�K]�N���O���tk�~��/�%U����iK�d����'K�"�w�����G*�{E�Rw���ъTQ؄���H�;x1mU�Z�L�
@��~$Z�zu`�ލp�����O�Ʒ�Ey޿�:m7;MH�{/�u��^��XD{Q�kz`0i���O�WWd�Q�E���X��Z��`��>��Ckd`�\����r;��Ko�D-	;[�"MO&#s@\�><>N���:Y����%Ɉԇ�R��|,�q˼n�E���FW��B}��M-`ʣc�x���{��0/��O��xh;���Z���Z��hΌ��n�M�) J����a
�7Y�����5���O;q6S�?,Q8sah	M?)ݗÇ-����xa:C�pys�I�Ֆk���@��վ@������&
0ZG�H*��th�N�Ƈݎ�v*:X1�u�`���S�W����Q����M���f���X+�IT�#<����^e����%Ođ�-m�Os���E-
y㴟�-i@���7�S��z[D�g�)ǕEU�������2 ���b�E����#P5 (l�ȴ2N�e
��M+ 
8ЯL#�S�I	<��9�x�v��Z���0�{�b�3�sN�]t
%��	)�����Wb�3������R��Z�}�����C�'�!�x�o�6�J^��_��0�w��!�J�
�D�.������-:�`,�S/z�.?^���ٴ�Y��FT��9Z��oԾ�L�k����jQ��(ۯ2�1~�99-�u�O��� ��˜6%�؁H��u6 �8���0�
��J#��h+�.;x��������	�4sI�4�R��?8�s?���yG�c�N�ǈ�Ht��.��5 �偍�E9��mhfFV$�^��*����	@�E�I a�N��s�-\R�'�6�nG>}���w���\�\ ����U3~cn ���e�+��t�ڈL'�޳���ߝ��%jyp�<���/M�\^(�-�n��|���h��-+����v�=�y���AQ2�#���d�
���?]����ٖ7�gZ�ҋ�w����͗���N�;������+�cߕ�*1t4��3bZ�9UK�,�}n���5cޝ~D�y�����-�q�{��^X�ٞQʘ�aQ)�.avQ��y��a����&�a"͑�J��"u��CgF(�c�v(�ʑ|EpΧ\MBD)�l%�[,v����q�a����������l'��<�wQ�s����F��W��J׽�($7E(R-�Q�B��j��H�*�A���R�Re��}�s�\�"h�}�>^��Z��x�r d�/�c5Kh`��|ƣa���˥���_�'�Ϡ"�g���.C��ʬjVr��ue9(-�+[���ns��u"f�u	NS�n������nD|ģ���V4�o�٣�h�+��K���$_:����Z���`��&�㷆{���ki� K��C���٦sQ�,�c6/��CF�lOi�&�l��;5@~s-=
��~��a�7�9��
	���[�������R,�?��c�l����r�i������n��]9�쇂X�r������p@|�ЯH�M�NK��q��k���0���5�|����X�'ΗW�-p����Ui@o[���y|��l��	�t�Z{Dyھ���=���F��r��I����)��~�HnB���,M+a����^��3��$VGy�s*�ۍ�s�er-PŁڔ���r�ˡ�(Eڞe�(y�e`W;���a�/���Z�a�)�w#����`T����r��#�7��'[0�d$���!\SHTf���b�X�u/{���kQBP���{�B4a{ऊC\��`m��$�[a�\�_��j���gЂ�D�(É��
�m�N�̉���\D�u�9P��RA������6/6��1�{��+As>��s`��8�g�Vaƪ��6�Ɔ��4�������uRRE?2E�76�ՅmI��ka��p�oU��9� W92�
��� �����2��j�ZNS\�f��6����v�	�A�T�+rb-?�̥��R�����l+$��phy�YS)G�X�uc ΂=�0�n[�<��t��ZO������]H��*��Q���^"3����H}�5qɚ��%����F���:�O�lF����^������<�o���J�d��,��I�z�Z� �u�^�cڞ�m��?s��+���K,��4�{� o^��ȏ?�"9E5�-"ٳ,�N�S�Y�����R	t��L��ѡ
�d��->�Q��:e;�n������ڐ��L��'�y��*̿3��j�A�*�\��j���83�����U��oUřM�p�ϨR�y����[^�[\5�	_7��	#�����z '�٩�-���05���X�� �_/��,�������]��GF���Zx�0p�����z)��Y�{�^�����4�/�S�y�x"x:��4"po2��V�@; ��3;!˶��g����w�Ν5�,�ԩ�&��vLOu�|��76;�b
;�����ڭTp�����#�;�J񩳎��>f��a�Ӌ� 
�%\�nZ�G@�+(����X���i9�cx|�7$Jo�6�"0���|�0�	�����;��%���=���T�t����X�bDW�qf�9�]|�b�?3X���n�s����K�X���s��Pu�o���&f���-J\�>?�~�o�����aV�� �����JnE�G�	f5����{vM��aJ���x
s�hn���3��R�k׃��b��Y���y�yc����u��U�eƟҞ<�7�Dd��m�L7��̣8���IwC-��I�d���F�Ns������-6��Z���Z�������F Gr�Q�S�J�ی�B�#3h��Ӂ��ޝ(��n
��4�6�=���#��Fy}�{�{-Q�+<A,Lr��Ԃi�Џ'������Dp��;|�]R���Mŗꖼ琱ӣ����޽��tNdRn����V�̢��m������Nr$��{������A�s��[�FA\�����m��T��2CqD{�]�5����"	˨c��� .�S��@�$��iP�7=���w$��"��L�����=�Hr'�c�u�5�Ɏ	'7PcCW@H֙t���	���/*�k5��c�θ�����˖�f����1���z� �s�iE��Im���pb�㩽�z��%��h5�ů�A����?�}��q;����=uh��"`�/�џ�]��ew\E�6wO� G�D�:�7���f?�r��P*l'�ᇄ}�>��f)���D�3�GY2�Oщ�Yqdql3ZE*��%A`#5D_��0ክM�)\v}� �Kj%%�}�X�!�A��m��EܭSR�նt��ޯ^�P^]�GS�Et��1��,6-��J�/5��O�_�X5��l�T�oO�n��7E�a�"��RX��%������� 
)v��#�i�M�A�KM�Ir��s�*_*����X�萭�8�)m�7�s��]~�%T?�ƶ������v��_���:&�E|`�������Ҏ�z����e�ʜ+�8�̷��L�p����^�w#ێȖ$B�!Ȅ�{W�s¿��4L:��/�1�ǫ�"ser����Z��tb0��1&°�5��)�A�%�i_:��b�o��4��E�����f��gG�W�qϔ)S"ط��Mز�B�q��S�U�>�Ru��~�͇�c:~3�/"tA�R���m���,*?դꡅ�K��:��0�)ƃ@j�.F����NN���=,�5\uQaڤ"�5���o�X���N�M�/5Ǫ1O�����.*�[:q�Ma2�֌� &���'�.NR�.	K��/\!�U�
�K�5om)H���^}����������f1������s�o2P�x?�Q��<�����SanF��H��A�5w���͚���9���[B�$1�Y(��p�";��z�h2?r1��Jbtz��U	�Fw< ���_�-�SX1��uc%N9.	8�c�t��4��dʴ��]��(jw��9i�����c̹>8����f]c�5�FdI�t�O �K3�I�A;˾�ղ�o�N�&fpƯ;�����X��?.vJן���H��D���<1b��x Aqy}Q�J&�&^���*�V��J��H��'ᶥ����d����Z�<����f�N�;�U{���"�����9��Un�+%6���>t���.�b�G�"���T�w�ƈ=�:�py͎����IT��f���]�[���mж'P(���B�A��U�F*�d�_���#�ڵI�#I�{Z�)lR������fw6��hY������&�u�Ff�����}i���οZ�/&U��b�Dus�;��I	�T�V¼^v赀�A��#��Lx���UƱn�hl(��\�ߚ�G���������ok/��K�!�|%����q�PN�7�*�K�<5À�_�U����8Lnv'���[5\\N����B����FxBg���D�O�	�a��R�R8�e1�eּ��KTV #����
kIV��1��#c8�VdxW�;ī�75����P����+Q��}%C�X�Ͽ	W_��;	�мT��
,t��F53�(mop_+�D�{�/x���_]�����|���ٟ���U�,"�	����4\M�{�J�k	h�u�.ä���\MO.��.��9�Z�M	���W�Oi���DM�FD\x� �VI��j�}k����-��R�t��8��D/J���(3��!����@T>�����Ч?;�� ��6����1î(B-jPrߛV��%Ѿ��_���q��m���f�ʚ���M����bz��)_�'%��c{����m+���5�ķ9����>�XPR�?+F��Ԫ7�"���⽿�Xj�G��L1 ���20h+�&�`�
�c�w�����"�A��Tm4��{�)��5�W�J�7�P�i�v t�&֛.�,s����������6�	��g�_��ט�}d�2��v�޳�e?�r%����z`���/qә%3Z͉��d�Z�#�k1�>��Ywx��=0߿�W[=�ao��p������Nt$�Cʏ��לs�}�R�,�4�QM:�l�&~_�5JƷʹ����͖�H�v̬�?y\�1�m�u3G���#��h �~9�7	�\��u*��P�:0��~�5Q�ժ�����]ڵi��˫�^������0L[@�J<�,Ժ]̓$/?��Ҫ�F��V�C���XQ^mFQ\�T0���-�J�8��z�?_��G����S�i��*Ь�U>q
��"���n�<�]9Z�>1�N�w�+�>#�d%��)'ڐ-���-�_�!u^;dpλ�����_�;�J������P��%=���k��3�'e�2V�N7$rd�t�ⅳ���H��%�7>��* ;ofD��'�ia��l��Kz�Ř�w�f�}����f���|�[Bh���:�������jV��/�@�����pE��iխ�O�,1�p��Dv۽]X��c��Ι���W,��F��a2T��F�d7�v�|71i���S8�5~������h�4dq4>ʉ�����%�N��g��i�.�M����C��\�"�T>�J̈́���K�;�	�����kKؽ�e�m�$Tw�]NYYJ� 6QH��'\c��/���k�9�\+�[��� zh���#�.���w��#lmUy%�L,r�яxM7#t�JſVI_K!�K����!k>=�H�_����P����me��!�x
�( ��|�5a0��"�j�߫4�c=��AA��?��X�If�}�x�5&�!Gя�8�2.Y]h�躾�T�+�_F��E��J�$�H��ǹ� /�ne/�>'��	u'K��}b��ѿ���V$�O¸��Dx���I����o$.��Jʏ�9�kt�O��&GJ���Y<L���@E����3�y����	��B���k�sf�4#�1��W��,9F���w.�S4j��no�'����߯�E,�L�=��y��M���L��[���j�M$����kfRx��keqf>	3���Q�������/\!_�Eo�a��Nx��6��q}�JD�8
a³�J���>�W�/3�R����#��RE��k�۬�k�A
ۡ�X嗑T�����CU&��=������q�j�x�,^�~v��OP&bW95�u�Xb�7>)�ϖK7V��d�||YC���=G��ٟ� 1����n
-�Pw�`i�c	�X%��u����|(�nϬO�,̈́���H��<V�Ҹ�k�W�7�]�U�Y��x��jp����"�~�)�K:9E�,:aB�� ��N9#j�Ǌ���?�p�&�}u7��S�`h�_r��DN;�*B�đ$L%�T���]5���o��Zњ�ɭsݫ� �z�C��Q��lh�ٹ+��KAĭ�� ��24�܇*�1:hK0U������'�N=�J�g�X=�&�M.�����ɘU��F��Q��L
�Cy�2h_���}p4�>�UZi�5�Y�q�^�m7S���Y�0���/I�_/pS�D�v*\斫�!;�'�d��[ۅ�,����#��r��k�������n�F�˚�s���/�k�J��B�1��C��І�xX$Ip<e��A������k�~�U�a�7�فޣ}E�"Aa2lb0�Z�K��5�J�&t��Ru����('0Y���2�H�m�H����o��ȢM]���/z�EW{f�|�K�����>gqX䠴�
�xj�T�2f��6���z�K�e/U9�쳠S�\m&O���SK�Õeq�mq���0dk%'�����d����{F��T5[PZ+��e�h�}����ߔsb!����`��?B�AtTX��%�m�?A{�M�!p�E���@�٭��j�~���U�Ȕ;��L�=/���q{Ǹ(�(��#m�~n��@��SkR��b*"`����(��D�}�ub0���ueS��=׷�Sҵu>	WXE{��%e�0QI�b�sh��Xݬa �G�[A��_Xh�x���6��j�t)߁����Ǆ���Yƶ�{��%f�۞v���(��!@��1zl0ER��2���{�
�8;um��:c����-Ejj*Gtuӂ�C�5�'��/q�x��i)g����-
!�⢚���gVCtq��kuBv�6MX���{���g����l+�zg\K�}E��1�.��|eA0�C�'Eu���K�� Bw�6�z��qc<��b$,��~ZI���k2�,�(~�Z<Te��*E�����@a�ys��`w;������G�LT��{�[Kl\�JGh�6M��;��@r�'Q�F���[�Ӌ����
W�O��	0ё��&҉a M�XuJ�[�&5��y��%��.<%^[Fw)ώ� ��B2۹�e^׃�&��-�2[��T'�}��ڐ5?��:��5�GZ�Μ� ��jo�_uN�ќ�?1�sV
h�3<3~���_������� ��KvB~-d��Ϟ���ou7jk���l��$(�� ��.4�����i�*��x�T�}]���AGuw�j*�!H� ���cCh�������~nO���^��*�8�����b*�{�Ux�~$<�Z�&�Q��F�e!3�*��UڡfGb�zMR��Hsd:\@��a��]��R���P+UV9�[��՜N~9u�tv��ծ�Sl�p�����u1^-[w� 1�AI�q��`���X��T�FT�촵]ߜ�֒B���Q�.�<Ơ�d����ȿ�Pˬ��Mq��U��s�UX��M7���������(�~���o3h��'�|SI
W�'�J�Xu5Pa�j����6[�Uf�< ������-f�s��9��;z�i���ATX�嘡�Kي��~�'�<�&dG�JĹ\�a�Dx�J���\QG	*'��-�	� J�䣄�?�����6Q�Nx�YJ��{ýl^5:c�n���Pzj�l~W�K۲{=���qp�E�������|��Q�xe<���_����;ZϢ�G��ְ�)�n�kr�gn��s�P[�����u��(��;预u���	��P�ʁ��/�3�W,-���5�=���|uB3�+L�;Ä�<�^�����o�j܋a_˪fH�(�?��c������!���%��ޡ�p��������7��(����2	\�f�4^?��cB��ǹ�ޫ2��`�/cv@Z×Ow�YV��K��' ;�.V�!�h�8�s�z�1q�? $m�#	axc��C%���[��jz������|X胁���$��y��d�/<D�f<�s)����]k��7g�[U�Kr�T���0��A�)�b�����ߗ�g4M*2 �Tx��/�wo��P���0|o�y���S(8��u�9��&�)�W.��r��v���N�)B������a��|@Ey8��z�).�b�XK �u���A�v�\L9"�:�\64:�/J�?����� i��"��i��A�Pf�E|���[g��u������V���z��߂:��n��2�}-��r�P�)�g�$=���.'�u��D�	��	ktN�(�'KV�)�GJ����컂�w���%s��Ow;X�Z��2,V�^֜a{3�`|�L|�x]�lwLl�[�g&��|�Fu�3�]��1Tߌ*�\�B�����cZyχY<�3����I����@���_��=a�,o��i��j��/�D��R�q�5?���p8.���7�bG+$�����$�BQ�`�܉��yb�"+�nk��\jȠ�	*G�\����G4����q���SiYIȠ�El���L�$���4?��v�9�W�u��d�oԶ�F&��I�	�F�V.��*uT_�"�4;�}K�7"� ��2�
*@7d��r���][ը�d��:������=�綬�N����b�I���E]ͯ#lR�b�%��|�r�]7����G�̶+�qy���qQw+w~ʸ��<`#��<�����������2�����%w��:�"�M�	<��dj�L�Z\��5�/Y9
�T��;ė&�$�qJ�E��� �SN������^�3���ٸ�sӘ!��
.im�b o[��yf�z��[<�|�����;�DM1F�pM�W2��n�m�\a�7�@x�HL4�l�@DE�6�!��#�t/YyM�
�������%�����/*��.�h��T%·�nqd��1�&�S�H������$ �%�o�"Ⱥ�,ok����{�D��8������yl�!cU �� 6;��s<~>��b���>��NZ*ҡp�E��*�Adt�n�O�!���ЃA~E,�kX1-�\ϼѕ�ܨ��:�~?*^.���{�9�/��M�챗�\����v�/� �4$�N�����8߉ϥq�HT����ŏn��Ɠ×b����X(BWf8��X\A����91G�H�7��J�z���I���pJu 
�W��@�n�R9�y���W�:��؞��̑"��1�ʍ����a"FP|���TW� T��������g��1֧T0��8�x�]~�Vu��u���[�b�����hb&q
Ô��mL���g	a=�%`˜X�������:�uֻ�9a��N9��/�}�-�A���(�lF�K+>*([?z�cv9��1ع]��΢����z=�7�rۺ��$%۫�Դ���(�N��Z4�pc��	Jy�w�Q�r9a���]�~�Z��	��zD>�O��ͮ{F�{�����π��o��6ȕ9#��^�����@G�ԷY~v9�a��e7dT�I��S"v���!���Q��y��jH�Z�������l��v<M���+����YiPV���.� c���兕5Cml���6�`�Ws���i��K��'�0?�rB�;�3�h�!��0����b)�f�_TuOx���zѽU��GBB4?��#x����W�1�@���K
/s)���:����X�����ނF'F�2��h����w�dT�I�0�E�˾�Fg��C(��2ϱ�ݢ�p�� ���$�C�ԲG�����|aF
�~[n���ڏ{�ͻ�Ϯ���qG��x�L�9KM?K���y+����,�/�;�%e�LN�h�n�y"�Oq�=Ƨ�;��g�a������4z�\0]=C���q�'��S�1l^�<̟���� �[�K5���ٸup��,,LZ�H���$?i�I�l�� ���N���F~3~,p�$6�����z�V�����'�S]�mO�E���I_�11ꝉ%�ப��)G��fm#L��ʢV�����d 5�C�mO1i�k#����UP����Ͻ�g��K��ROM�~&�d��.�eJ��ʨiM�Ĺ|4P��&�X]��d���x � ���θ)auJ(��O�l�;r�`���s�0>�[Jv
����쌳`W��F���tK4ǝ�孠֝}*V����p{�D2/ñ�*6�^D �9h�)iMg�;@P\���4��1����J���:�eރ���qЏ8����qo41#�Iv���踌�JN3]z��/�;1r���-�D���
 t涊(ʻ̤uKa0���*�,D�)����n^L��r*�H1�-�d�	j�`Ǹ�mU�у?�z#���ݟñQ�"h�!fRt�M� �Nc"�E�#��aU/�UϘ�����m�[���@o��w��vXx������=����H��	�[<��+2��3Y��n��F���w�w+�,�:�Q�n�$�Vs���L&�㢸r�0�K������)��$*�<��l�Ј��)��OHHҞ�tc�%���ѢK W�� �3��ꘝ���� 7���a�qg�xDx��O�#jn' �7����H��ݖ�I����qw��b������	�s��e�$�G�*O |%�.��q_� �M��n��<�f�0#�{ۄ��;���;����������i�i7��uT<�Rf�{�P9�5>T���+��Ȃ�`�tI����U�0�0�-���7�	0J�#�(5 �{�.��6i��3K��D̊�#-ZL�N+k���S���YGWЈS!]���Enކh�������~�4���4�� ~'�
3�19�/}w�bB����F��8l�����_�*'A�y�	��R���UH����"�Y�{O�����v���F�l��;��v�ӥe����J�,�Ny)�홆����ȕ"��e���6K%)r"��(T��Uy�RB�B�ȁ��c�]���2�@�lQl��٨�t��|N��\��=�ЉF��+ǐ��s/�D��#L(wu��v���Wbہ]�`���	�~�9ԇR�˞ �N�4�8G�#h~Ɨj�<���S�߆�!�2@d����!o�̫d,P��ʫ�m�>�M�&��u�Śo����{�z���^V��N��F�P68w|���>�TX���c����m{]RG���T,����
[�`�ߙm��$�f i�S֛��|s�Ȝ� Q��^V����r���H.[�f��W�E8�3ŀ8��4?F��?f����U��:��>,8�4e��h|��Y��=�G|���vv�2Vk����g���!���L��n$~t�^�m�����e����`K��6�ɵ4!)KФ�Ae�>�i/G���l_��\GT��c"R)Ų��۰�*�'K�����n(l�A�ӷ�܃�HM�� "`��rO8Ǩ�7�dإ�|⬨2���X��<�4��dtU�{�](į��C�'�E�F�w]~8������%0q�+R܌�֨Y�ÏU#SH��?MC�O�U�!%�}��ː�ќR��;Ǹ���-`�eS�+4l���?{�[F,_[]�R�8L��xJ�M��� �<���*����v�����y��cǲ<D�Jq^�nsk�h^4�Ty�cZ��u�M?{�E�\G��W�����4�>&y��LoN�A�+�WXV6��ƚ�D�b��g�g��H��gS���,��u�?6�U���M�8-K����:�Oa�<���0M���BǏ�1�aڻLA6���9	�;ꙧ��������JVG��J��Th�"T�Q�`|����'�49b������p۲W
�Т�(�;�R=���p0@[�*C6�l,�T0�iVҌ��������,=����eA�_J�)��ͧ$�㔋�05��y���J?���+�PN�D�`��%�o��:�v�9��bT�:��w4̲Q-�J�I �0(C{BR�56s�w�2��g��<@��ק�X�7�3h���7�m�x?DS���_*M�1_�E��te�����Qˈ~��ˣ}�2�ѷt��fx�Mt�6��;��SGe���� ,0��*�X�㊪�*��O�N�`�kL������Y���B�צC���t�u۩S�H�ɑ�o<i�#h�v6c1A){J�����(�>����@R�y�F.����t�*�ï7�g�����ɝjINxi���qnȖ�}+��w"���9��#S�i���ё?~���F;GU�@�>��_ם�|� �r�鲁�ݩZ����>�k�N�o����KC���P�R?I�z�\NbG����ٿ��Q���z��t<
z��d�C$���DF��q3I�~|��+�v�LR��o/��N]� �Cq�Q�$ZH1���4�˵H�@��qyQ�QL�����(�S�X��Z=�y��F�VԧL�����P7➤��������"�^��J5��g��c�
�8M�
Yަ�G�?��Q��;c�����!o.�/�'to��H{q���C�"��l�4k;c��i!�/D����W]`���'�Td���b�I�!x�� `_tC�ه�M*�c$�_wFn��9,K6׮��:xzwӈ�0S��9FtE�|w\P�I^&=�Q�)8�Y������f�F{nu���i�J�ī�3�:�Uk�T����\z��D�V��\lN��^*����+�5d�5�k�FE�����:vT}tdB(M4���k�=��,f.��ڿ����~yA�	ٙ��&�Ja�S��i�`^�����b��{�T+2{T�}2ϩck�\+B��Nw�7vD�M�HB��^�v|�{ڈ���n:�,�Z��^U�j@l��?����=r5�@+���p�*�_�)��!i������ ����Q�,�3��[$K%̯�EDI �K=b�e��ұ��NY�Dr� ��i����d���WFyB%�6T�!p��BQ˱�8cs!��%�%L΁���Z��9p5!�8�����23�H;�ǐiY��Ԭ��(����qP�ͱH*�����I�^(��}:��{��0��Y�	S��9�K~C�A�d(J��C�ר����Am%R�C�._��l�f)�F����v��V0�ۂXD�ҏw"y���Fo��l��Bd�Y�=���_�n�i�z�6S��� �K�Vw#��w@]���C�$�u<��w:�=��<g+��:���gFkom��}!%�t^�u��gƿ��T�|4-�OY���'�Ɗ�3�ҞT�$4X��U�$��C�9b��^3�'%j&N�4�ԋ�t�i������\��[��'��gQ9,��v��@:��ڏ��"�I�޶.���of�a�'`��n��[ӝ�D�n���8#C�wj��l�y��E�|�Oje��F�3�>�^f��@��)!�^x� .��iua	��9��X����| ��ͶH�l9_]Q��_��`�Ҝf���e�Ԗx�N�P%*��i���Ĺ:7i'l���k���d����b?�����=ݵ �gO��:����o�8�W�ceς���4*/J��=b�׶��BxI�*L���gpr�l0t�+��6�y�~,�-�to�aMb7���ke�v��9�L���[.�+Xn,�vǳ��w&-������H��iT��++�H�<�-o���I]M���=�f�NM�1����J��k\c[5ց-���x8Ƕv�sV���Sh��38J2Ow:+x��#њ�T�eW;�yJ�l��<,���W[���C���v�Z�jjѷt��|�8������F��b��<�]C��XboL�J|V4��`�ZΞ�}�i��|̿v��a��B���� H�8���8C�>��Gq�Ƿ1:�S`�Ӿ���_�d�a��ˮ�goU&Ϥk���B:��wWa"J�
"TӘ=�������U�z�j�a�&�O�5ﱕ�r0*)�YL��Ҳi�X�Tx�vJp03D����ׅ���X��������4=|"���D�&$�G��������Ix��ވ��'Z�~��F��S�T�%>%�-ur��K$�{��9�;��ӄY���t+������r��H_ʥ��o��&U��%Kd��b~� �NT�C���O|��������)v�����j����/u������@m3����;�b�S��������!��=b���o
��o[�����l�/�(�k��p-�NM�*���2W�)�|��Y�!����`��j��s&z�Y�sTc�\��(V��h�C������˱OL]8��HI ̬�u��wh�#X�"�N湮��x?uU.Ѽ�����e�����u����0���s�6;����	c?�#J��g� �Q����4�ʐ߫_��V���jbM��=�hrsa���:�T)��qcE����zv��d� ���(Pd�ֈv��yW����E���;G�;A�D�QPٸ�-�^��e��t���<�6J��ܔ�@>y2I���؎Ğ����A3�r��8$�f��`F W�6^q`;�2�� �{��¯��S��H��O��33#g$���ƃo��/�!L�آ)BI_]I{
ܔT�h��J<�U��J֍o����F��]��tځGK%�^��Ϻ��һ*-F��􌝼~���
�h���T���)��}�L:�u��c���#�)ے��g�2��,ItVR(�:�&I\0O�i[y���PIw���@8�̕�Ǭ��>V��K���XY�a}���Kd�e}��jro&it�4,��8U_j緛t�F����9��r����t�2��]�#�m��Vҭ@���m��g]�N��U�����׊��'��BL�������С������ �6pJ��?������T02H�mp_�
�6)��2g�Ͻ�v�`k'��/������f���?;��K��	g��6{B����kh�?Y����h���\0y�2�%�ĺa�RQ�b�eŏ)$b��J�R��h~F�nq޹E�$���WBn�𥤶Ώ��NGT�c����6�����7$��f��q�x&x�[<H`OA� D������l@ѿs�PG��G����Z᪲FN���J�H����$�}��Wǎ����e������ .�IS�O*� �b��	NI3.��>*K����?��q�3��0s�:��A`�s]Os��nè
�+h=#�#��>���A�UY��lV�/;���<�����`����{a�dx�XA3��}H�Vg��A�<�"k��K��9��|+xM.�������
x:�Ⴆ����s?F&�n���K%�����[��4���������k	�i�����nOX�:nut���?���84��c=��3�)F����5nn�gkN���:vU��p�hZH��Zt�H�e���l��gh�4�E��f�
U؇_!��WvFyj������u>��ԫ,��%��%:d�����2�*�2)e�[dM��KD����JH�M��g�.�	���/��
&�9����i��|{X(�Lu%g�˘��K��b����ӭ��-��XZ�(؋%C���1�?O�<�=��n�.�!�%�)��9���\�,o`�yw_%EE8W2|ZJ�h�s�h[aY#�q�{�9�S&��w���o�:���J��L�2�tz��� n��J��w&|����.$��k�SG!l��0��P=�{�aĿ	<Sy(y����.g��lTA�Q<�Kܜ��뭕�6)�;iH�Z��i�����0K#��W�
��궙���hm句n��̀��:��Tp�����G��_��X���+�f����3��z#S5	�p�U�c�w��W�m��KQ�	�C#3�Y�G��&Z�3��g�#TH��X���QY"���d��b[U"+{z�M�BΕ�u�6���/����ݧ��A�4�¹n�;|2�mBMG�3���S�7�1�JϮ�o���� 3��f� [��z�c�l��u+��"�gmz^���K�jM*��y�]�=[_��}�1W�0�R�;)�������b�L�f�@@�Jg�tp��4�����7�����!^�7��Z5�/�,�,�F{釯0��J�g��L�mWr�V�U)9I��ؔ�'��R��� �:�w}F�"+�&ׄA�u<�l�b-ک�=����Ɉe��®l-�+ъ�1�3�����S;�"�<s�	/��#T�;�p�z�*Wc��ܨ���ƪs%?U%�D%@ ���F����x�8���f��W����4��W�=3�������!�	�LK�XɈ�p|��9��`��|��b����]�"��,������4��^�������[�]K����Jkm�5�X����r�qp��y2�ak,�i���1P2!�-�	�A�Z*�ʝ�s��(��������^�ۃ«k�(b\�|����!��t� �s,]�fzP)��4�F�m1�R,���oo	�K�|^��>B��Ӳno*R��{���c�W]�]'S��c���2�Gh8͝�6�+�;���/�KC���Y$w&^Y�Ŝ!z\ˍ��β�0�1��f���#����(W�Y��L��I��M�������u�� ����VTs��,e"y�`��8���Ο�e��C�0���ߪ�wTÀ`���˹M_���N�L�9�Wy\�ݳ4���{>TI0��n*����T)V�?6��32���V��7�:5	�H �HX����W�5�~�|�GUO�������@��Cx�ʰ�GI
Nm�$|U��3������;ᑺ�c;�B��T";�&��J�$1�������*܉����
��53N��
�Bڬy�t9t�d�H~��;���� ��amt���Lr� gԀ����w8�`>�M�U��_���=m�#q�~��Q�D��po�5x��������e5|(#V�Dw�/�F�M�ƪ^���1s���~�}!r�dg����PT�ԝP)Ѳ�t����y�WL^����鎖�Q!PS��2��_pmf3N\3��F����M���ٹ�c�? G�����7c�v���n�˱J=˰P�S=�p����4���8P���3���0�3��p�}/� h��{�+Q�s���6C{g�@����H��l�k�V�������\���GF<�7��s����G �� B�H(l���k�!�ORl��q�sGT*Knd�`<L�'�e��(���+p��Zh�(��[�U�G�X?|`��G4�'B�)Wj���|�0��S'��~��}ն����Ul^���9V�<��*��6�C�`�!.x�S<�X[P$WoG���S��|n��o�C�V�/9��剶�g�y�p��}��𕢔���Y�R"�v���^����̍S�F�
� �q�;�p��(�yV��
�L�C.�2�s�� �o~�����cK��;�#���ߘ�c��E7��n'��>�P{�{��4���*N���q%����S���NBfqA5���9�"rCX�X���ʃ��8��00ۻ����a��ͺB����kj��h$/�RF>���3�q���@��T��VK_�pc����=�L�˕y]�.瞾�c�J�t�-B�;Q�Rl4�p�q��E�3{���n`�?j�f�g+-��(�H�3�f=�t=��!�Εxl:G����%���S熜��=y3�̧�G�y�hw�FRVu��~���v?����������V�� l����ߘ�Kk�VS0�����t�@Kj�p+0A�B�P�K�0�rᎺx2��N/��QW����;�8=*�3��Y�t��=%c��pw�ԍa6�)�)ni�a"��n)�\aF���Vq�����oc��R+�^�q������G?e�C����2,�l��gN?�̀-�=nV����v�Az���R�8� ��?�o�Gab������v�o�)g�1�{YF�))�b,b*�u�Q ku��
T�.d�rg�y��i�)��V՞ h����V��k����܂�Ҏ��.,4��Oͭ %Dn���ſZ���y@ o�m#��$��j�t8r������W�j:�w2	��컥�P,��08f�ډ����h>;�\�a��W0�6�C��������k��}�\����������+�q�����8f����9
�h�Yų���ڱ�_�T�\L(��e0H{T �����XX�
K��G���I���e�7A�f�-ÞFy�:3l%�[tf&\�fh3�#���1�7�梷ˤ�[曽��I��'-���������[�@D�=A���u���v��s���	j��@�y@~���"�tV��'�Y��B�:^y��v��̗��O��X�6!|��m�w9�	-���';�Q�ԩT1E����Kf�dp�n8��G��$ؔ��t-��^7���}�M�T,FEE͆�$�~fU9���
ܭ~r�ZQĲ\{̕r����N�ǁJ���ݘ��̑R��d��0.yϽ�ח���A-D튠�Mb�|Ûv��G��\c糷�<��W���.{�?���"���������4�x��+DV�`�f�m2?-A"��|Hb�5x����7�M4��o���c,��(BK�i���l C�XQ�2�m�뢝�) �^M���Î�ʦ,�/8c)ϳs�K�<c�"��O��?< ٪��mo��'�D���K]�m���hd�sO�L��U	J��v~M��N@Cڼu��x�_�K�ǲiH$BoKi�Rsv��E`�`q���!�Ѧ�OC~�J�u
�Gf4<�.��8��0P��pk��Kb~�s�7ߞ�Q�P ����|�?܃z��{y���"B�c���3#-k���^���R��!��14��/�ş��R*6��3,��{�m���,Wd��LNK�:eM�93�zF~�4�����;�9b�굟�zr�Smz�E���p� '�3� ����K��� *��+ݤ���:6y�lϪ$��K��LO��9ɎG���\����(����^�.K�V�����rZ$,z[�����_�_ƿ�&�Ex�W2�|PX{�K�{�B��lo��e��"��=���G<�bF\�h�D�"\VW�&����5��W��xd<4-}��z�S��30����O,<5_�R��D�_���:yy^��Ւ0��F��D%_N�%\;�����ˠ��8r�b��r�F�*gvL(�Sҧ����e�4�Ǿ���Q�g�\1ΛbQ3;Aa$�Fa�@*�K�9DT����q��<z=N���Wj��"6R���E�Z�u�Sf��_�EwC�7��AЙ���^
�pUJ�E4��YId��f�oG	Q���(f��d���W#m����49Nfg{��.�&�^�3��k�2�q�!z��͚;?@1��a�T\ԙ�w��{;��9TT�a)�o@]}�i��߽��&1��*W����}�H� >`���M~�ѷ,ك��9Q[�z���x���?;�)**�8�9�p�Fp���	����]��4����y]Ћ=$�OQ�g-�Tu&��;!a��4*_c����ŚC����.�ԯ�|��g��d�eR9�řd��:ۡV���kI�ʃ��_[�EZ��\Y�6�LP< �ޞyg�aԪ�Qo��!�VX��k6�5՞g��=��,������G��m=aATUI*ş�EÚ�?���I���3"]�&Z�/�/�UBkϢP��(�n��@���;U����H�uf�1-w��;�1İf^�<�h�/#ҋc�ڭ���Á Wĝ�=(;S+g_�EGh�Z�[Z?�M#A������������Q�C��.[��k����]�)��?[�p�o�Ț8���GD�+;騷�\�u�}��g��lq^��=$��$ڶ%
�?�k�߷Z��lek����)+�0>�*y�~*�������l�o#W>c�W�������a>X`��_$f��"�� YI;MPrI#����aXT�D�G�d��p�l���t������� �f֖\V���@w�f(A����]\`���e�#��N&g��ǽ�y��w�A��\�<zO�Շ<�/�Ȏ�} f�zZ�mY�Κ��Fl��;� �~��8�SZ3�:�Q�͌�_�{������W�^��l[�,�Ñ_k�`���	ac:s��3�j�"��(1k�v!���c,�;���4הC�*h'c�ţ�='@�b �i�}�$�<�G�oz���/���b�/&h���<٠a��/M^�ܸ��%
X�$�Ì�<��5�l`(�F�C�x��th	���i/��|����	�I����P*�������:4a�4�܃�7:7�ԣUJK/�E��`�U��}��!:��:CR�o��Ί{\��XzX�a��k����+)�Dρ�ō�.����_(�����d�d9�tŞK״��\6
@����lW��٭S�ǢlS�d:k*>^�]�qS�L<���&���<k�L1����}�V21�4*a���S�V��*�4�(�l�P���9*�3ȗk�v���������.o9�B��n`[��	�ص���Ӽr���HX=�w!e1� �:��p���)#M��&��O-dm~�Ҙx� �X"��r-�G�μL��"�����n�GQ=�&���Ц�kd�ήR/�X��e�Wo[^G�x�U�U+xRt)�g���fGE��8k�$���I�v2�B&f徆����$����*���(�x�`Y
�7b$s�	���6@1��Ùڹ�*b����^C�ƨ�b���LC���@�j^�t��o�,�U����zU���l�����t���0�o��M��9���o�U�g*v�@���b��3���l'���i��L$^d�� �����,�I�0��jk>�N��w�T�L�p$��kDٚ�z�+��M"��y����5��F%��%0���k?w������63�]��K�R}����w�4�G��&ʨj�@uZ�/n�x�����!��Y*{�Ǌ����X�Ő�ئ^�*�_>aO�y��=���3�(^��b����)-��ym;��vM;�ǖ�[~�|�Y��O��z����,���c�!��b�����4&���_�!m?�U�/�G?���U�mD/� ��+�^°����4��Uy(k�d�e+(릍�<I��h�/2���T�yŏ�YB��,�����g��68��z��J�)D���k�:�/C$ƍ�^�Io�h��W��FAln�\͖Z�յe�Ɬ��������C�8C�*?��[O
�D��l�&�u���\۰*�]}LTV�hH�(}��VE�Zu㪝[^�7�'��2-�Jpb�С�6?}�z���^���Eˡz��}�*�������NdI����V$��m�q �|x|�@w)�����NE��a�3	�p�GɎs��O?�؛�K�sib��U��$� � ƚ�gw$�/��0�=���r�.!x�O�#�����K/F�$9�����7M�<��EZ�<S'�D��X�����5��#v�1&O�w{�˷S�.A�cO�f*�����a\ �w��9ӦM�~�;���3!�)?W�ك����5]-R-V��8��`J��(VsP;3���y�B��@�_#�i�C$����8�8]��ek��rޘ��M%R�W��?
�>��߁���2�'�&Y��o��X�����nG�ǎO��0h����o9"��䢥�:,�Jef�3�4̆���3�Led������j�b|E^=���r>9�R{]=A����`�x��.�mL{w��nx����9�s��������֪���J~f�z����m��i��;gc���z�]ș�-'���A�_�6($�䕤�?Gy���;"��ܿ��N33����{��4�b�(`}����xG�f���~
:D�%`;Դ2���Av�1���ի�Q���YL��2)N؀Bn&΀�AF�MT:�&|�e�<V��03�,A�Y��˭^�ZL�H�)�"��r��ӵ"E}�mY f:t��	="#�@ތɛ��3D>w0�L�lg{ծ�o3�||���o�M�|�ڃ�,�����%n��E���8���_[!�",J�ݤ�� �S"A�C��m���W�<q�9��Z���1é�)��D���\i�꿌{�_rW_�w+Ut�e|���P%�(�|G����U�)���֝���AF ub�˝[��5z ts I?џ(J4Qv/���=�U���@	�5H��>Ag`������P���7��H�@I����ާ�媚��f(L�K�X���B�O¼K ��V�~���$Ϡ�86M�EN
ݎ�˻���e~">���n�rX��H���r��0��~�����xƯ�����&R+42�����g��`�.	���̎�������t-���Y�3%��&[d��7�u���ZQ��# ���N'!A�\�'6��^2���~�*8��G����If���91� 8Q;���{R#�9P�tF	w��T�d�zؒSA&����I�}��#���L76Y�u����	����K�/�j{S�H�:���H��X #�d���+i/H
�pG>�[U����W�j���)���Щ-��YQ�E�pGE�ěz�2{n3OG�b�j�� ��x�z
h��f��v���Y/�H
&���&����I<�J�FmR���*������^WG G��na��~�Wq���\�0���s��|CO��� ά�����H��[�Dݭv�²&SLi���p�l��6�1�%Xc�q�iJ�u���s=��FN���qw��iӠ.����i�:��>��I�2�I�C�@�C?������Ǒ��!Ii�j��ʛ.i�ʸ%�� %|���8 ,�:����Ai�S{���Eo�)nTR���	Ƈ�>�mǨ��D��\�'�����מ,�M�P�Wꚗ�2�Ҝ���沇���M{�̾�J9�jӞ��Q�^�ݕ�>$�n�b"�YƐ֑�pg���`��.�ٳ��rxKt�}m�VqD�O�C�1��Y�$�|��j� �֪lҢ�O����i:Ȍ�4����m� �9�;!�.���k��pB��ؚ���?���d�~��z�>�qW>��L�o��E�M\���R�����xU>,�V~����4�͘���N�"(���͡D���{녨��~X�ȭK��{F�<t�O�r��c��GD�!��b'%X�`���_�I|6m���t�d� �X>���>R7��}^��
�Z�q�׆���]�����̷<a ���[�"b�����}�՟O��0���(awy�(�����=]`V��S�����9"�W�}�>:w�h� k:�w�:v)W�6�݈ԕI,���#X7%j����~$�W�0cU��3��O���}a�<]��l�媢}����L�F"$���7^(�ά����U���F����D��Ч�};BN���d��լ+��_�dQ�؀%׸��9Bڱ��3�!Y]p��8�z�*�v����4X(zXH�3�禩]�a�tpY4S�B���i���F��Y�g�y{`Ƀ���ŷ�H�iw>�T��'�|�HE͆�F�&~�� ����~�˷I`�2�CP����x��ƶ�a��e�ޔ�Z����K�"�S�Q�WD4�s��v~f�r;�WM��y;��J|�獑Ƙ׉L]���q1���	��`Y�$@�f�~\�m�%��0	B��Te�Sڽ�^�������A�6#�[��V��$��ar�u�%��\�g�ܷ�BK � *�ł ��P��@����� YP�6'�~�=�v�sM�Sg��@�F�d��H�$�|x9o��_�=�KP��T�����$c��R��&ǣ	z��B��tŨN}��[
R�6�åj�����w��P`�����n�	�J=IM�ڢ˟�n����o�����n|��M���D�8���r�f+1�qd��;�L�՛a�7�괌�`U$�Q��+���_#f�1ʎrXfY�PқG�F���t��p�'��uM	M��<Z �5|?��zIZ��oE��W�w���fBځo�W��IΩI���$p�Z@�zQ��� �=�����������}d�l�ܮ)r�"�h����2�,G�M��0���K �{=�i�D�7�[�����=�;���[M��9Z�J����3S`����J<���T�]��Њ;ŇT�!�ڜ#a�A������$���+G��u��n9����e�i�ga�'�b���|��,��r#G��r�fSe�� ��Ȁ���u	����s�"ߨ�y�%�e�������4:�����i1�����M�{g�ygY|F��h0,��%R�5����%��@��	��CYN:C4�d��틡��*r���� �L������J@�d6�.���<֗��~6�l��rm�$��g����}C��!
z���K��O��w�%���|���Th^e��Lbc�5�t��=�/A<L�f�R�GO��k�������`K�:�e*<���Z+��O�}�Թ&O=F��T}fNY�!��	��Zg�g3�h#:?�R�lj�8l�y7�Hq�Ҁ��y�D���/��|���SЀ�P�P��#�D�N�>��I���8��Hdǀ�q�8AN�L��Dp�ޖY{����]|�شާ��O��ׅ��G���-a+9%�4��m~��lq�
��CW^T�T�۟r�Ϙ�Aǫ��=�ҌQ�3��5��6,����/-������Ёs^�pi"����4�݉��:�=�@'�?�*ly����h�����G�l_��I��u.)G��0H���3�>T����>��\dR����&�[1!&fB�&U��A�rL:7�F�`
���4��(59K��ڨԬ�,}��e�^��!���K.�$U�d�<5e1T� �ܼX�0IP-�5G�m�ѕ��	���ր��C�MI���C�������c+/s�|��i�I.*�?��V�������	A��7%�I�{�E���7�3"�@ZE�W��y|�+x��r�ȉ����j�Y�1Q��H�W,y&���S� �2q;8E��#�!&}9��P��-
�k�.�#˪�y@*��s��jL�]U�t�x���,� �'�K^�|V� #/f��Yv[�g2�L93j�91��#M
Qc��ϡmś�;-��qJXv>c?n�y
i�jVG��Y��������8��أ3���֔u^]��N�x�w*���<{,l���U|)�j��֒B���������J{:���Y���sa��<�Xiy*����h�T+MZ�n|i��iP��ny~�Z�L�8دŗZuD2*�����7E�2;����u4�<�=Sb���zݫ  R�E�w���HP��0e���A�����!�Vuh����ʕ���2 zڑ���n�hc��Ֆa��~���~]��Pį��� ���/ ��E�\�2#�z����`ms�V) 'O��Ҩ�"՜������ 2笃���9�ș�E?���锟! �v�uW87��<k�z��Ue����M%�����fu�8��>a�{\��XE-��3Cb#&��M�J������%�{ .���k��s'r/u��j��C/�z��c椈^��V���ɣ|� �PS�WU ��b���n�h�Q��dt!>ZR?k�wp���� ��MS��G
pp(-�Q7��H�N���Q���l)p�QuQ��	�r�'4;� �VD^`������0��9�-X	��<%rZ��	�����.x�J62E9�ܪ-���� ����~¤dI�
�@gs�a�wK�~d�BQ-k%̝5`Z�����mĬ�)~�ƣwE,�]W*��B�LC�1iM��1��>).���J�Hk]D%_�5��&7������	��2mR��ynr2���r��Ya��a��W��)�.EٞӖ���/ E��W�2m3Y%·(�v5�O�Hk�f73�YU�{��5:�CjE���<1F�h c���1�'�$kCy�b�[ Yۢm�eSC�嬬����~p`�aV97q��+ė��I���Ѳ|�:@�����!Z�����
͛f"�Fk����5�������<�����^�[�z�Y�)�q��Z9i����� !Lħ��{�R���K={���8��!.uԾ��6��ʓ̇U9∡7;���̅M?��3#�D�]P��j���������8vm��錰�h"gz��в2���������:���\�l�O�&p&Ъơ��}Zi���8�|gf���U�׊8*���r~#���!i���OYr!H{s
��k�xA��NzTq�l@��%;��.Q�Um���^��n��v�B3��F�@<�<�u��#s��-������y90�+���W��M+�#=�%)��
q�f��0�����k�t�re0�ʤ{Ƣ�n�C�0���3����aJ�7�ش-���G?�,�P���9c�A	Y������ս0i}ro�h�ԯ�4�ZF8rwr��D�d�u�S��^�Qe���e�_p=��0�����l�	�oٔ�P)g��A�a�u�9$�6��o�RR�1�~e�F/爉ܧ��J	+�繯9	\d�w��9*`�loC;��	�@���.��kqH]h�}0ӣ��O�����&`�˪pSK\��I
�����Xj-*;��%R��K��Ñ4+v����FMEd��X�&0f�U�]-�o��-����BD,7�F�� ��%kܑ"�di�����[p���y�k{��	�m���Ok���+-�����Y%-�ʢ�&�Tf�z��2kAꋮUz�*�2ڔ�i��ƨ���}�0@���r�Z���0��P���(2��<��$q��^�(vV�_LfKvT��;���gi\���@����E<�;�􋊄I��p�̝���+����.->%�{'$�Dk������xoP�^�?@��E���˛Ѓ4�s���Q��H�ȡ����&ck�l�l}�U|i��ۃ�I�s���FB+p��M��$%������->�G�̯1����l����6�&��+�ܝZ�`�:T�$���.���+��ܜ��s0;��	�X�GJಹb��[�:�Y��R�Ҽ@�jR�-{Z�Bڥ���4��؆���{{��צ���j쭙�I�G�	Ġ�^�R��g6ͬ� IO�+���3f3� �^5ZB����q��z���,�{jX�j�ʁ�_�'�1�����źW�	଄���	�a���'8�y���@�W+U��lX!ڰ���AQq��+C}%�=�C�����ƨh�wm�<ɟ�C���	�� ��H���m��o��ۯ�-�{"E����ݎ0�Ӗ��1Z������U��I�Aʷ��r��˕��d	emo��ħ�i]$X���(�h�-7ӄ�	���?��^rΒU[�k����:��<��yQ��G�˰i\=XJ�H�3:f����f+M�B�p�I>n��}��Z޾+�V�}���<m�Ҩ��<o����x���0�[�˘����^ѳ�aQ�s���xgT��2=/���L��pǓ8K�	�g���iӒ���ӭ���W�G��.�H���&���t���g#�K�Om�[X�ãUc�ْ������L~n��ZS�Œ;Ī��kĴK�������c�~W�����@��B��²��$2�E9��Lt��cF*�O�1^E�1ߣ��l�8�I6cK����
�1�@�@�?g�jb�vֶg�O��F��s.1$���k�<�E�_�L��H�(;t!�\�Xm� �z9CL�䋓	˰K����� ��q^�HYݢ�a�äʁgeD.o@�A��Dd$*����#����2�*uo#����H��E�g�aľ� s ��E6U���YRE1�����o��\�n���Y^�Ů�01|ġ���@ ���x9�\<ǇQ1��f�#��L�P�W�;
�����9��b̹�k;�D�.;��zn����ٳ�� V )Ik@��	H�췖� ��{5��T��i%�����PY.O��4y�cU6[d��+��F����"���^�\����K���"t�g:�Y�%y�j�4���k�\BTք`[q�W��K��)��9(�.]ۋ|��mP�i���y�4K�+�?) b���u�){>�I��D�����d��=/]�~.x-����ME3�X���d��^�qv�}D��۟-/�2������C�i%l�"�&#_r�u*FO���cu00hE;	�Q��d��O�t8e?�������:\ƬrC!�4�gʒ<",�����t<� 꼭,��XMׅ��rb�0޶&ɯ��}����3d�J���1���J�����[%t`���zK��;�ȼ/���t�eKo�%����kj����]�stz@��=+ D"+����<_T�>V4��z��HV�.���ǳ�y=�i�2��]�M:�)pYk�ڻ�D�����c��k|��^<v���̴đUA	C��y�d����l������N�(|IK3���6�d�����ZP/r�l%��<W���ӏ%�SU!p�`&�����ؠMT�ɮ�R�2�$�k�ao�O��.^n4!|��F���'N�#m(B����զ�NUcW�6�%`����)���F����65w�d�@�o���&�ț?�]���/Rj�L/��*11��Wru��h���-p�˥�H�@�E�lW�����v
�q��Y��D2��z��뫃x�Fg%�yBt���p��º/�b�6������(>P��uW*W���	���Y��:������3�R1*���-���"<�K�a���Ò;�����ȡ��
n~>P��I46����:�W�fh*9Y	T�	4�Kߤ�?��
	�@#dx����o�ͻ.i�H��W?�+�)�4%�F�U^���Q*&d��k��/��)�(_@�K�ʽ�d�(��It�y����ԝ\��~ꁣ�_ˋ<���5"�����jF�k��9:��F�n��ܜ�ov�p����������]�� G6�%��h. ��k@����w�ʳSBʢ�i�۸c�KA|P��aj��_7P��<�eR	��-�p��npe��24y�T�	��������ۄ��WB�ۗ�D�>�8eg��?�
a�Q�mFk�b�ah�]�>� �^��2��$׳�hШ���k��l���КVF�7*���-S=�C����Q8^:�|�uD��Y�P `!�x�f��;.��>��EG��@���f25>K����������̢K1���4��ߡ/�����;���Xˉ�`t*'�^�rg%�%<�G\�K�d��lC<7q��N�,0��eC���;�n�k{x�X�;�LM��*:ʮ$j��A>�`jc4�O`6��Ŀ-⛣&�N�h�0P��V�BݪM�ަŕғ���W�Ir�o���ߵ�"x��Л+�%�%�J"I�c��F��K�7�!l�zc��3�Wf�v�:F}�y�[��%�2�<�7�ZZ1:��7�Ja��,]��Wm׬�x�N_,\��a< ��VA����2�9�f¤�O��{���:~�\gɺ����E�0<�!zK���0�4?�cp0��b���^�9��)�hWN�.��F��.��?Y�,4V� �V�iO+xR��*M�\�#>��n��Wb��X�I>��)v�V 'Y\�d�pg��B)����l�AS�$'����$�9�BG��ʘ�{��i@��� ���@M��Pt	�Hs����
c�����4w�N���3E��oFk5uzt�q��ӕѷ6K8tH��p��0�`N��=%fc�����2F�([B��S�~3���& ��p��l�f��[�FG���*B�/D��b(&��Ҹ
դ�*��)��NںR�}�;d�NĪ����궉˺`�B��W�;��p����l����rO���q4��Х�x�_���<c�	DN��,�ڻ;�OJ��i\Y�W����-M�q$&"h#���[�A�j���X�>0���X��Bj�z7	=x���T�|�`�I���Ѫ�����1�5��Prr����� {ܠ� F`0լ�Z
�Hx�Y���7��1���ޚ��e9�z�z�7�Bu#;���8X��2���aKl�����I(��jd���1t��Ú�A��	�?Yn�)~i���lre��_^�����gee�*��ML�̀EҲ��xDͫZIq:�� �զ�rU@�G^��y��ݡ;����l�Od	;�φ��]`���S�2Sd�OV\����ӊEp��B�G�o%�������K�"1X��B���z#�F�7I/R9l.�N|^ �oJ֮<,ѩ]��F0߲�(L�,ER�� �ؼ��\�֨������r''F��浽��q���#��)/?�'�E����+h$+O���co]YN6����+4�̓���F��%7���0�M�x�E�#b�"e��fOp��Lb��Q.�װ��GcN���J^�w7�rG�������hztc�����t"�r���,G�ҒG�I��M>�?BA��J��P<���i��P�m��\)���d�X�~���t�?O�;��@gj-��3�����Lۡ���1� �+f����H�����X��5(��,��l?NBE��M����z6�jS���wojd��N�a~t�m���*��v�x�F6aX�b����6�8Q�&)(�Z�?Wl�
.%Q�>�a��{RT�2 ���pDs���^�����/�9u?��'_���KF�E�
ڱ"X��f�b|�S�1����עCg���5�� ��6�x�q��
�q(Ҥ1�w�oI��V*+�|.۳�����==X�C؇vlSۍ��U�F�WB:F)]Cg���tN瓦�'D͛�w��l!Y
R`m���@�OIc<(���x�4F�-ʦ[8�D����\����*��|��
!��K�k	0ٞ�K���g������J+Ȫ&D����kQi=?�?&�F�F:m�<��B�v��]���(+�j٢΀�(����[��3Մ�ccZ�iv�.e5��"�PϘ��������IR5�nh"R�zQ$]Z6x�Ӵ�@/�*=��Nv?��H�z�zx*��f��^w oX�����~��|^�:��V��5%p�\�&���*�3^���P�X����FؿS*�[§LL�Ma|GGq�厲v�f!�˧6Gg��xG U��+e�$�ED���n��5,l�i���{��*����G���r�Q�E��'� �R�_�`Ia�3/�"������讛��a��ʌ�BOW��ք]���:���[%x%I5�&�yˆN+()"~�ڶP���rz[�aZ�Y*�bC�^�-d.��0���L�J���x��v���_�!{�oX�b���R��x�+��8.��N�{�ib�/_�R��OI�i�,������ �H��E^(�Q���X�׍Q�a!���,u��q裄��Z{�~'�����q�`����FRf� k��?�������� �#D��+cƸ�q�L:�`l��!��\[�D����r����y����C�Eڍ���7C�>lo��ބNd�wB՗Î��~�"��"������Kctg�.���ש���Pܵ�� �\�=MT1�kDD&'$���G�qjd@h�%p�<�����m8=����쪆��9�uu5��2�]g�4v����2����S�8�w��%ŕ�V���~f��Nv��A��C#�d�I7��b`�7��T����Q"���P���������O���m��^����b!�'�5�6Wd&�����,L@���!�l:y�]�Z��v��A������pf>?>��5����鷸��9.���7����Kޣ�Zl�R��p�Z���n^U{������<�,%��4qŧ`������Ew��⿝�����]��'z�/o�dk��7HK|8/�r)���9 I-ޟ��;蹘���L ����J���
Zl�JT���T�������F�ǭ��D�H�ן�kuP��z�_�¹`w��̏�c���y�VD����gc�#c.��~pJ�������k��f:z?��:V���>K\�ը&7�Q�BLkGd�mp�j{0��Z��X��?���%���fi�NN�U��̚{����-1uރq���x�vr�Η ��.������ӶSoDq�r�Vg}� J��YW[�*�O���1�j���([઀�b�6.�z�d}ԇ�}?Mer3R�"�'U*YK`q�tבo���f��<b&��o�Ȧ��x�e0���*~�XJ� �yv��ϣ����Q>o_�{�v�(��'���wD]>[d<��T���mEBձ� ��8~U�{�<�v�SlȄ#��r�j�s�p�,|}��?�����5�\p0���0K�X�s���xm�<����
�v�um�A�ő+�y�U���E�/�^�u�J�ΰWٖN��C��w%�G�X3���Yi�m�,6�<�]ҁ\g��ۍ[���Z�B��i�Ui����b���hɞ9��ѰV��Ro~��W=J�,9���< �V�$��|oD�Ļ�̮��)d�(�˖��ײ��䖐@�K�EZ� �Aa@���$�
j���/VɄ�ٶ�y�\ھ����g�-|6T!f���/ĿAq�h_>n7�*��r�Tߤ��%w�c�����+<��z���I�s�PQ����[B�9ɗ�_�H�Xk�?T���1�BL���os�7'եْ0��`���^G?�����.s��w��zT�����T�3��.	ovh�nx �ez�C���z����k�Br�̶f5��+�:!0�Q�&fI"��'��ޞ�ј^t��'�ce� e���l�l�Ճ�P�u �n���~�M4��¯~�*�>�];�{�t����R�a�NV�����ȍ�a��0e��������Fі	�,�+n�YL����e�L�NDc+�> s�l�Ja��#�ߵ�KTx~��7���6S����\eX��][�:ꬓ�=疉�A�ӭ�����
���o����b���T��V�:��\�s�~K���¾�*�~���w$�t����B��#���P��� �����l���罟P$V�H�!��OP�v�;�����ݸ�dj$�0ޢ�|����_��\�5�U�Oő�#XN�/���֨;ѐ��>"|�h�
w�=}���Ia��k�<|w�gA>Ji�r$���V�^�v�#2r���8����/(W5�M����d+�FWA�>ފĽ�q����VаZ��.���bY:���
��xI����æw�
�͂�����[)���t[>*�k�J�?T� ϶�Y}p\�L/Q���p(����|&_4�z�$(�&y}E�t���,�z�g���b��8C�~��B�?�U�0��~��y�	�>��|����gD��	���a��l�T�m�\"��"(��n�Xvff�:̪�/��O�Ƽ�t�T�4�A�Օ�M6���ߔ�<���ڷ�j>��g���'g��~����V������i]��f*-m7y3u������L���y�+�CR�#6�P�Rk�Ȟ<�yX7��NK}�o��~Z��S�;NŇ�|���RW(��"��u�����i2�[���$�J�S&c�؞N�����Y�H�h	��E��W������I#X�ոS�Ly�����0���س��"Q5�x[��|1��s�Ӿ�m��/��Қ�[�������C��`����yFnI;��n�'�Ҏe*Ir�O�� 0gN���"i���s^�d+2m0��4ȉ�I�Ϟ&��آ�%>����Xf�@��,��N)�(4�JflM�x-*�G�|�~�@����ZV)g�{D����$��p:�Zѵ,�� ���a.��E������[9W����dJ��_��q����Z7�Su���q�V�g&�SQ�%9��%�\�uhL6�w=X��`���r��L%��|����a�d�������ۅ�� �A]������mOY���Ӧj+��4~�����F�O�=nKE��,��	�l�!��Ѯ1C���ZfmD␆5-<Kߝ>��_e�B%iWa�n���I��sh����~�����H�Ti.�E����m�V����U�tE\s���f��o��"��@���у�=�k����FO�/��ZԾHk�٘Ug?m=4ȩ�+��)�E@D3�9R�.��7)1��	6�l��+v�o ���O�d����"H΃2_y]�D�4h��C��q�3���R���/T>��aI��b�o21�	xg�@�JіQ-i�R^M�h1�i\0N��>�8]3�5(Sؔ=�+�qӧ�,e�*��B"��˃��Y1��(SG-�K�
-��8��no�; �.�q:>�|��/��/J��.ҡ�}�.a��T08��Wi%F�btYx/
IU�쌄�QQ�/���))��ᘓ �w��
N�8F\@�|�~5X5�a��d��t��<9`��4K���	SϘ挡v{l�Fv}�2U�R�����TK�c�$�S��z�Jsq�@W��MH�-�]���wwnA��r��Sn��-T�͕��a���l��ZB��L�9lQ��d�X9D���2����9�2vE�E�>㙬�)0���W�P��glk�9j��O�)�Y�}�f��9L��k���:b�(- 8xݭ���{�{��B�	4['������]nx�ߪ�S�\C�4dp	����ZP���4	�__�Nc����a�$�/4G��)/(�ɬ`݂]�����_�L�����v�F.��	�I-�Ϋ�ѱG�K���7���u�켨Kl��$��U����UB�徂ّ�1Q�L_w~�<�,J�wW)����{����E}�]�}�9Ʌ�0���Q��
�¿������������yD
�gI�����t 0L��3����Ķ�Ga�F��mF'�
�&���~��d���ۓ��o�\r���.�V����U�����W, ��/�G����|��M�Eǈ��w)
[�����_W;�z�$;mf������ =Afj��G��<��k��G!��Ku���.�t|Ð��������T�"f�{ui��2��9�hь3���,<R�ч�Eh��8;����f_�Ĭ�T^�b�y��h_��N7�rݧ����G�h��	j��������k�@@hF?{��j���d����E6����w1�/_�REd�F�>;��y�:&bD�ah����^Z�jl�:~��.A�?Ԙ���s���Onq����J2�Ԃ���>ۑ �"����V�EEp[����N��=��CsP[c��%��Z�1Y�Rё>,m�(�f���]��aK< �ھ\p�(��yf��y��Y�R<�I�\<cd
彀}�T��(P�l��S��H���s9��-5�XK[�n:s�!�L����k���"ӝ�?s�C�r�p�o.��!�gB'�cSq���$r���M��L�4���X�&q1�㐄L0n{�{q��W:�� �Q�`�
~��.�p�W˥1�h�Y�`���G��oU�/(W��ս��1��Ί�y�8 R͓�+��_�0 l��89���:b��/�����T-��D�
�Q��
���6���7�ĂYc'�U �世<�s>�u)a(�m0{m��ř-��jRS�1�,�*���Q?&p׼�AA�~��a�U��٣�C����R'{m]{,ǭ`9o�	��R:����+���Bs"uq����6D�-�آ���1���W� x� �y5�l�1���+ӏk��y�J��ްM@�+>��`�\%�m�fq{[�j������jC�O&�ߎ6V.�=��%���0rH~E��ꡡG����4�#�)��Y�����E�Y�:�=Ȩl�i�΢n� �ϋ�ʎ[�N7�,�[%�K��> I������?�$MS�gx�"����T�|p��U�onɐ�dAk�.^����E��;��ꭣ��2�8CR7����E���]�q��s�"j�0U�JX�:�[�]M��Q0�� ��x[��Nu��1�HJ��~~�nM� ���f	S���.K��3s��L����3<k)5��ȗE�Q��Z�7�9z�ݛ$b\c��wJ!�����岜�:���p=ǊCUjU;����i���~�HX�.��� Z�U�D:����
�X�1/�WrD̾�e+��}����m��Pr�� ����.�4[}�qv|i�qԚ;�C^k�~����lתYE�TG&���F�o�~n�c��[ ��tF�(D��I|ȭo��+���r�8�xj+���[�&��Y�l/Ќ\b�I��q��*�;��G������K������g&N��\��7M.�~��a}������o����7#5��s�8^�<B� ����������`(��*�(A�2s���@v�޻(4ɠZ��{�폕fW��j��^�Ҝ���ޝ}��ٵ H��B��9P��Wy��_2���ߊ�Er��^��$��9-�md���It[0�"F�l���'v�N�jSY�dy�x'��<Z/���C)i��/RD�����!�����kq��q�m�r'����ZsG0��-Bلħ���e#�N��t�ST�JxqT�Gw�<�<���l*}!��R�6J��)�n����9JI�'�Q���skb_�Z.�\5J��ܻ�󗯛��x��9�^�O`�`+ol^��<E�f�e�q��6N��6����l�t$nU�]}+/��J.D��gѕ{�����H1Cj�9W/��KU��azD��/�^�|PY��䦵���`���( �ӠXuίgkd�M�12���(2E��8��d|��ԙ���`*��8�����K�������W]���(�>�G��k�rJ{J��ʂ �ltg��U�Q]j�"������<�Sf ����n9������'�f���b�Iٝ����V.��"^Ym��I�i��K��R�:�]5�3�9�Q�t�I���S��!�!b��n.�eyV�����)�ܹ�V� �c�q��p��(��z�_��ߋ�t�j�1��t��\����յ�V��b�b��0ʮx���z8T��YU�r�ڄIV�*�T�	�ÍY��iAyc��(CS3a!�E�2�W���WR�|���MS���`�ܓ��ܚ��<��~�ɡUH�����Oπ��!�8Ϩ"�P��P ��x}$W���R-��Qls��ȃR(&c������^7��ٿ��d=A��d`A1(��5tAF:^�p��Sd`���tUI��ĵ�����K׈�-M�6��ˣ��)�׺ @C8j��e	��L"�.��=m���s��,��s��<V~�o����)o@��} �4[�p'\!Z���%`�&f�w|����:�Næy�}�#�̏�@w,�����1]��פUZؚD�a���ea��R��`�vN@���֟�}���q�?űV1��@���- ���Ҹ�U��7K\�$)s)u�s��O0�{YD�؇0&�ǫVN�<�w7�:��Ʈ�nt#��8^�d���]q�iY��S@Hݸ�׽h��y��5d�Ꮔ�� !�[�o�ڇY,���]�<����X�d��٭�����eǟ7��nZ�N1@��M��B�͚��L��2G>�3Q�t���S	ٚ�84#`�ȥ��;�9Y�� ����#̋JGi>J�q�7v~�]¨���1�UN����p�pP*���_WfS�oAs��o���ʦ�\8"��e�;�~��6�*��Ur$�-������A��_΀!�]�Ui֮�2�/c@n@�����T	[�`�A�N��i�U��y C=��ʸ����G5gsMd�1��U��ة�>�&!�,��B�k�^�[t���V��kC�Z�|�"�y ��JxC���d��|�v3���vs��=���_`�_���̦rح��\R�>F{I����RiXC�j����4���<�ЎMUr�X�K[m�*0����d�/c�;6����{�\������WG�s9V\vyv�a��ݗ.�ïT\��w�"v��\�|�hi�S+y0��1���ÎWW)���/�թ�W���
�qz�+�q2�ag��Ej��gһDKpV�pl�_-
�ِ�����A�K�[ 4���U.P2���:�@C��Z�؊7���TQ��]E�t������a� ���n���]��4�ټ�^ ���o�6e�@o�sT�-��1Ȓ�g��t��n��\��k�(GAYw2�I~9�z��0k�d�!j=���a���!,#p��kv1#���Hr�/r���^'�� p���/u�p��3��5oU�5��i�N���u��@Y��YSQ�<%v��"�
:NR��u$�2mG*z#ß���x��8�Y�ſ�}����.D27�H�4�o����TG7���͌�˂ڝ����1Xy�.n�3'w���O8Oj�;4/F]�W������%�ɔ߷�����t����\�@�j�vM8ǂq��<H��yb"-ga��c(f��Sj����Ԙ�����ld5/;��$�h����,E�І�V�������aZ��i�_�<W?���nv.	o{m�ĭ�Ѹ��&�._i�6 ���r_z�ߪC
�M��9B�^���+젵����w�`�u�&�f�Cw��� ���e�����+�]�W� �1������dqi
W 
�G|�0�m>%e�) �<=8?�i3Os����.$/d&xE�FԐ�?]�4 ��2n��	{�Z�16?U�� �q�v6+���ҽ�Z7t�_ո���PS8�Q�r��!Rj10�9� ����Q�����ײ15��x�E�@��e�+=��9��f�9jP��>��4K��.7 HW�	�\B͟P;�g��_NU�/�mk�cD�6�e�Wzde�8'�����;��I܅�Joz-JN*uzH�����J�C�B�½�?/�*�ZQ�4u�W��S� ��=bk�����~���F���<���0{87�Ôy[�S��;9�UKN՗mVH	�7����Q����N�6��n�o���smJ�j�h&��pQ>,O��	�w��ķD� x�?�׈�/����r,Ƞ�C4�]+�8Z �?��=�ì�8�9E�<m#�J��<B`����'��ؿo	J���/����͊�#,t�M��G�r[��i�ɇ���/O��z ��ב�Ձ�dtz�㨿��O�o�[ �t��|u	�
�+1o��r��d����lE�3�1���+E�W�M�υ�%��y����")��7�u8_l�_��2���]�)�f��IU�`�Air��{� �օ�M ���=kv�x8:�_QK�4���Lv�Q2j��;#�nmYVe�j�����i�c��
����������l���b}�NK5irᅍ��F�cl�[����C�;�(3C�������_ÒIОlO����d���q�Ɛ�h�G̻�˧}Qw�G���/��|8�[���1�3���梿�Be_h`��B{���ҫ��&,�;,�Ef �9TA��/[�{�z���,�h	�Z���l�qN%��<���SKi#O!�fn#ApU�O����ط�����7&0G��0���e�+���P��y��;��p������l�o	h�ra��H�o���s�������k^��_�e#��B1E 
���� Vk��ېU��(nxv���ԟ�I�e�Fѐ[L^U���Ţ%��)E�s�3��[��W.�l�wV<2e'��Jp@�Z���9�u,��D�$�R]>P�9��}�V������d�?���zC��`O�e(&V����Y?��M����>Z�03��ӵq����&B�ӥx��Rz8$�9Ō�!Q-�T��!�c6J�d���P�j���sY�+�.pА�L��M��)�5�'�\An^5I��IDۡB���k)�7X�=�[�]�B '��2�k�Də U�Ց�^a�&T�'��,���NU��N"����t/:d-��E�-8�a�`I&{K������5f����sdx5U�����^�D|��H��%G?8"<q��fu��x�ݠlh�(BLq�eB �S�ea�P�ef��L������>��q�:y%�L�/ݶ�Ȓ���� V��F������^�'J�"ۦ�G��7u�����Oo�h�^���ޑ�-��oQǠ��Л�B��d4����1i��"�~4�}]M'�J&֡ګ�h-rڝ�����F ������%����!s`9�sh�y��Z�suL1��oT*Ez�T�S�
L>5/��Y?�Cf�n��߳�z�F�Dw �[3�����h3�C;�0m�}���SL�~E�!�T1�`��!�/g���Y��i>��a�s&HC�,4*�!�*-�B��J�A��C�C����=Y[	�'����ʻ`��&��J'�oϣ;���Xm;�*'xX�-Y�b�¤��D�z�Zu������������s�`^���S�W�5�S����"&>yX�j�m (��:V������s�i�lwi�W�V�q�� ����]�Yro���r0�57d��@$�?��V>��0��1~|O��'-�^��{�O�JE4:;�������.�?��?���:G�瑱�w,��N `��%'�E��o}�-o�ҳX�?�9-��A��m�P�T�k�Y�w�-p��ne���X�	����ʳ���]�8#9+4�8L5W����ob���=�),@$bqe�� �c�՝C3��n��c��rm��P�_��P�Z_�n�a_2�e=��T�1���$sF;Y@�U���)��n>�/(�ɪ�����7ѳ�78��|���ͫ133�/���!��RߗCj���~��u�3���;_�a�
X7�J\4o3�o�����%ݘ<Im/5�#�t��,2ˤ;�.,����厅��P��d��{?q|��8�/�B�0<	�����6���
�s�pI	��{�l���_��E���K��P���P���N�PXt�}@�J󇍯�(��e9�5]^h����~���s��8�8�ax��Bv)�<T�"n�=ǭB�O�% ��&�b!��pM��>���W��U���mՉ��T��iW��(-�X� ���i�΢�y<�P�yv�Q��=��<�&���B b��W��G<�b���ϑ`Ä� d\f�	���LĹg:N�VS|��!�@~]���p�)8�>{6e�"QO 9Eu������cH����Fk�����a �l���ZIS�Y[[L?���Q���@����u��4�V��UE}��~-�8/jWl�oE���uW��8;��O_�S��u�M���^}��(\�!�6?�񚧎��B�����^�mS%�e�]����������<ބ��_�#5�Z����rn���<�6l_Eu�.�0\n)���?�.���D�����$���k�^U�8�A�(D��P��Ե
-�YT��~�>IM�Q�:�0�	F`�f�v��d�!�
@�SX��o��+H� ka�P��k�����?<!by\fQ��>V��T��=0���o�������Z r����++�$�<m�Cʅ�b�����+
9}=좋���Q�(�'�q���W��6}�,Xi�R#N������}�1<}�A�/�Ej��XY��E�a��{�?]qcu��i����������n������^����4m��<��߲��u�T(��U���{�H5�C
$|iW�~v�M��C�����U�L�bA��3[$#7���$:�ߴ���+������Z;�o�X�r���"��Wɢ۩�еFIX���B �2R~wH#�s�ta�_^�{���cT.�A��4�]�6����Fe��"�W���J��Ĩ�Z�)�͒r~�fs�_4�$|�n<��a'R���\7�W{Ɂ��4)����
��*�`��2�]���
:`c�tw�r�H��2�/��֝g��z�Z�N@��������%T�J��M���wH��=������m#.����U���n> ���z���N��W�����!��ب��gBK�9�lp M�]��d����IT4@�؆m�����k�3C��}�Sv"0'h�̚��Mk�J���ig�`|�y!�b���Ţ��,kT7�_Q3��=���R����ؑ�&"�]k�ݠ�o�?�%!QB��Ny�5��ӄ�f�U����[���D(�^2P��n�V���W�a*b�e|�Ry*/�!���H>��_ �8qʵ&e��m6ɸ��cԎ����pΦ�~�y��},��v�.J����\w�Xc]:N ̹����9���q��a����S�/�{u&<!��k�
�{>]$,*����?����Kx��|j'�ğ�Z��[D�Ǣo���p�_��w�W��������^�<�#Kf�E� T!���?G��St�Uhyw@�җ��Э��>��WQdQvb�����\�>18oZ��i��-k�Rr�xɆ�w�~��a�~�Uz3����pY&���d�b�w!D�՚��&�l]I,���k��qW�D\�=�f�85c;��/��e��Σ?.U���"� ֹ�5v����%i�8=����	���]Ѝ-�~X����w|�3���'���T�0.F�?]N�C8����?J\_�r�G.?�Ak�V����&
��A<��C-��h92���`{G$=��vl���I`e0S-Ǐ�Q���B
-������̓!,�!ȓ�pu�d��߈����4z��w�}<�������wcF�6�}-���!�d���>�k�+:*���/ڋ�,&�� +ܜW�)�V%|�Ø�c2��H{��@E��2�҇Ao&����
�+��=(�8�[������|W�Z_G���*=h�~�d
���(kW�y4�0 �0'�7*ʠv�8V�u�t��LRܣԱ���c2l��pS�VB�4h���a`t>�9��bٗ]�z�EsC(+z.�t��r�SA�M+�$R6q����u�a��E��0�R0,b�����t �lhw��Z�>5,�L��\.��}�f��k��#?GLu�Ё�D"��9 sE���B0����Q����XxYp��=	���1�i����(3���`��GP���O!��5�bl"
wnc���?����\<��(fqw���h)�(9h��Ȍv'&���dR��]&�z��v]�q��3h���Zr����S��I�v��߾J1MI�z]y�ʦ#��N"���7<��W�IŤ;�m�$i�~8��@�c�Q��"�n���c�K�biؼ��,��g�hA9��5
�=�N�a�I�j�ԑמҐ���3�U�:J��H��xj&�Ϙ>9g��̟o � R;�[(Ő�]7�|Ҏ�l���)tG�*D7�j*��4� ̚�egU�f����o2�ss�����:n��ТN:z�دA�����5�G#O���;�G(Ick9���ש����")��K�.�sn��)���Qj�g��|�p�l�%���2���MJ6i٢���뭸�m��h�8ÁD��O�I�!��i<�\�⎀c̤�y�\qF%QW�'��f���N�/�Ri�׏����q'�Cf�V��^�rb�1��*������e�����t�Β`~����1�n��b����[���:^]WJ�Ҩ���8P�3Y��1H;�ͪ�Ec���,D֛�BN�!�C�)u�ɱB�v���^*6-{���x�ٷ�<�r/3E�q�;H�.r�� 9qfc,�4���)�	EW�|��;L۰'>��A��1&��S)�MT.��!���l�eX����R�'�9��+�<@�Y��ްFŽlɾ^�q=g�pn������ѯ/z,!��y)�C�s/"{E��F����b5���Z{��ޭ��)�w����uk����TM�Sy���@⦧���C�b.�����8+�~��J�)|lF�X�w�ؼ|�ЯmF�OU3�	�a?=�'p�$�� $�#̭���9|��P����O\]3v�%�����% Fo��<�d�_1��I��|��Yd�|�(�K�F�VMB�5;7Ԩ!	փ�UH$>V_u���/�u�j���x�<��+%3'��j�J*��]����Z���l<�i�i�CHo3�+|Y֏�1vH�@�@,�g[rk,�mSʇ��; ���u�k���c׽Z�(&����X�7�uG�L=W��J�m�RB{�:��b%�����c[	/�D$!B�d��G�@z�؞���e����J)ꌲ��;��_�K���σ��-�kX��T�3�㢲5������ р�t)�N	��#�A���w7,1��G��i��^�V��V�!S�LP%�c`�Ϝ��<�T�v���k����3�m+��Gw�aF�F8�pJ1�!����8��o�y����̆�<Y�v��s��$�Ţ�P,���㬷*�&e��(�3�+s��~����q!�e��SD��,�$X�B�a5Jj����.��ݶ��6�3�j����!3¾%?ʋ��:~Z���$
g�0|ʠf�ώ4�X�N�]Zp֘���Z�i'Kd2�\��!.r�AS:3jU �i2Ө����'�6F`��U������>�U�$g�����d�%f�HX�0�h�&��9�����5_���"�m;w�T�1h�V�#����@h�X���@�Pa�x�զ�Y�C��M*�lG�Ǳ���=�����)��[x4��W����X-)�$b)�o��I�4Ltʰ��-(����Π��~�����u}�5�������hȪJ/m�t�<��n�ΪMۤ6࿗��@uCB����RZd~�WS�u�u�{�~�Y¾�<�u|���^������&���0d�:���VY�����$����;�Q<f(.�9ǣR\��vq�����F�V����-E�Ȏ�Y6ǫpk�����D�;��28�4��o���&���-�[��wRza@�i�b"	�x���ѐw_/,�#� �uG$|��~�k'���~�����55t*����	:��Q&�� ��n��<E�kꞌ��U��;�ͦ{l�CD�6c��ew`���U�'2G
3�	�����_��sSY8G*b>�`
>��� �}D���/8� 0���%�_R��S�^]-1�-R�=��_���4n<�`��QL�v��Ivx�q�(�b�B��<qA�,�>�q��b{D�c��oFr��"�x��D�󖠀QrJ�:�r���N�@��:+��L�'������姃�p]k7ŵ�qz���|yU�0���ث�@�~�NK�T����A�����P���p��7���̱�:�j9|��c��d���$IT{/���2��$��V�TP�>'��*AsY��/�>��H,����ekN��v�LML�I'��{�>��Q�$��&���ߗkx�jL�ۄ\��6WNb�()*e�`A�;4?�-�ӺؒS�}V�0Wǜ�]�C��z�-�4�+.�\o��A�l/�j�� �=�$� �'=l*��QQ��r.�����u�kl����}��y	9�c���z�����@'dAA��Gh5Cֵ��>̳�0�Ei��=�@�ÍЇxWS:�p�ᔫ��{#���Dw76����o���T���t.R/����6�A��~ �2��IAȝ;�?zL�~�������[�8�o^��Q�K��Zx�e�����Ⱦ�tB
4� ��lK��R�cQf�N�ҺϽϽ �4�@�N����z�T�e���?�v��s��<�8�����· ��(�M/�W�L5z��Ҿ@e�d�� ?�����xq8�d�a�$D���˟%�a��^����Ѵ2|�>@﨡���x.�s��W��>��x�q���B���B�8�	�;�<u ��r\W���2Sg�な�|:<�J�|�$�ēr<A(��ITٺ��4s(Ȼ}>t�p���N��l�N���c{��7�l��� ,���y ��g���d�ؓ��ԼcL�#k�S�P��d��)ƗM�ڲ�ό��5�ǄJ��%�rJ:{��N��!��fi��
p�����R	aq����ZR�B�(�z�@]Sh���Gy�m`�we.U��t�u)�^��P?p�]��ZC�e�>�E���_h�EJA�ǭkC�9�p���P�,�\�ᔉ^�A|�h��D�b�-�<QB��q.\R�o���M��4�3���v�'��""C�S��:ϊ��W�^E�W�9Z�)ݾhH-�._�"�5w2�*V���@�"� [�?~i
 �|`�+�`(�'���.4:�����V�dm?�_�w�C�P�H)fۚ�kV�����Z-�LV���4ؤ�ޭwXh�B/�uʭ�E��֫ �(n�t�&��%�]�!�Sj|%z��,������;��O����G��X�0���Z]5�$X;R��Jp	�m�%�*2����Թ--��X�g���cn6���6�+M��h*a��"��4'�l�vC��n�1G	>:���	:����F�岲�=%��J�s�GJB-��Y�G��& xY91�U
��$v��:ͯM�k8����ͳfi�6k���*f8�G`\�ez�Qr�e{Z��'�8�B�έ�-甆�_cV��d�MV� ���W���ƿ/�B��@yH�(Z�3��N':� �9H���d�x3g
�3�>����O�����<p�kW�%�KDW�;���|�mQ��O}�\�?��a�妥c8����*J�9���q	�MX�$�rVciM9hr3�����E��
(���Ԃz`��V��l�y�,}��[���բѺ*x��+��ND�:�����-�z~��bi�z*o|4���x�=uɱ2��+c&�X����_������`amP10�ݨΙ�a�����.�A-�d}�{Z�ys�O�k����z��8���謌���H�@f&R��q�.��r�~�6b]Y_�}�rT.H�-���+��~���ϋ^K�r��ق`����Xx����L�������v7���\��Fa���[�l�YD~^��6�5���!9GYȉ���sN�8��:����z���"��q	��ay5�p��e��n;F���Qg�=���#@Ӆ3�7�V��u	4*z�8��j[
�tgm#nT`���^T�b=>���&�Z�?C�ӫ�F�q�f����Gt��|�>;J���l�ܛv̟rȠ'l�wP��z�%�U~~��}+AVc����@?n��+���:or �/akK��>�d��K��3ߎ�CJC�~�T�����%El�I�܁�G�q�:"� �򸏠��ȡŻ�lv$��O��q��+#RG5�U���1r	��um5��7{��Ec��)���lL޸6 �a��[�	Y3���G�M�W���%�5<�W�k٠��ǂ���R��glGT�gY�Ɩ�пk�7IJ��ʥ�H��#ٻܿ���ᴍ{��>����~�:S�šxp��������ْ�Hs�y��C���٫���7Pn�0��L�+����{�؟c_���6�~��ƌ =���������[��kBVc���g%$'ζr�1���>g�q�7�m_Q��:yN7J��W�����[g��4���rP��an��ōho�M�xǙ�o��{��bۏ�'�_����|W�R{���Ec�����[�Ń>�Y����ge���v�[=��Ur�܍~L�Go,��K���o����M�$�"����9���������}�k��$U�Ѹ��ɸYB�r.t 1�|��9pf�bϩ�RYf%��c� �w3�[26R�^�sɏ~p��Q�k��#(�Ԉ������ֿ��셡�Eq�Z��#��&x��i�*n�{��Ӊ���c����c�����:��]�D
��ݗ�PiĞX��o_�'�@k}U�3��`]�[Ά&+^%5T�1����[�����R�HW+��Rv�+
�Ԩ�^�H�TEx-��L�Nս�Y�Iڎ��\�qL�Ή��!C�=��D���=���5��9����3a�����00}YW(�T E6�_��ÿ'��oj��kd����i �!5�Ƿ�S�hz��t�P*J&X
l	������f���G���g˗�t�W/	؁�҈[
�Q҆	Cp'�A�aMC�	�I(om��h�a`	���������X�EW��𨌡��EL�M�`��6�m4�[�P-��B�}W) V��5��p<Y�6�K��Z[�sT}*4�%��N�.W�%s`��<{O���6y��
0SX�ܳ���esN4N�>���U!�Y����o��� �7{������-8�ӕ
��W`���T2�K�3U� �9Ο�~!������k�f?6PH��J4R_%4I��.F�	��rN�������]c��&�"�%�3?�2X��ȖF�>#���c�g��4�;���ώ�S0�Ŵ���N��Q��2l�"Y�Smu��P-�=5�u+��}�򔲙
�;�ؾ���=u�_#,vYUƑ:��j(륡a���5y��#j��)~"F!��5��>Q�x!CI�Qp7��\�Y�:|�f��<B��e���VX*|���1�/Z&br4i��q�.��V�6<
b0�^`��N��n������Y��0�P?��8j+���j^�K��ԕ�������;���_�\b�	v21��_r���0�����r�~X\�E�z�$�t���9��
[X��0��˹������}J������{��Aڸ�C�蛔y�&��.�����"�Nn�߾�R2J�E�� ����	k��J���F��5Y)P靧�+ y�<x��V�:j�Gh4=l#oStO�f�Ć L�I��Z�q�b�?9��V)����#��W��)C��.���w�ya`%t؉�URl��!N@+Y/��u~�E��\ ���*�<g��U�ff(���	��/�	CW�?RBjƳ�%���5����D��-���}���fNO�z�d��j)�EY��m�n�-Ʃ��wƢ�{����hT�1��"Oi��Y�Rk���N�ݿ�Xpd���A�:AH.��d��!&�C���#�;�gr3"M��]Y�%�@ �Ѧ7d
��W�gL�0��_�I��4��>�r��e�<WG	>d�2$��#E_>r�X���kw�N۰�~��+|�ur��=qO�H��˨8FL�5�m}��l��	W�ݾ1fmH��5�SC�݉��Ů��ɟb���*�P��T�[�hR�;�
��;/���K�������:���k_y�����V��F^���������M?ȣ�y��DH\���:Z:L���C�E�����.J",�;Y$7��Ɵ�����D%�4h� �Ҙ��[ ��n��;1�,z�+2��JM2�)`�}��;�G��2�Ҳ��ֳ�k{��K��rv|�'���*>�n��n��˒��I�3��>�k��B3h[s9V;a���	e9��&�.^L4N݌��>�ѱy(���9��nn��D>=ع�7E��(��z�@F+���ߴ?��lV.䒐�N��}��Yyy��w7=�Zޘ��co��{C����B�P��o�ר��Y�i(��:���ϗ�ي���	��M�}���AA��M�h��[ꊏ�����7 ��K5�~����k�K������o� x`��!��z��~@�c��߀[ ވ��5,����o*��G��m�outy���@񘭁q E�D��ʘ�s�0 ɑ�a9{��s"�=��9+���a=e���P�4�!jn�t�� �/Z�ԥ�ۡ��P=�P�-� �|E�>o+.��7�41j�M*�zq��1I��<QIn�|���]Ғ��C�:{*#�.\�������Ű��̩:&3U��l�N������6��Ʌs�U�<`�ט�J�����ݻ6-g�Jw��%�$b��A��=3�Q\q��hˇb���Dӑ@;w_�{�%i�=ax��'�qk[�2	����|�T��V���1(�.մ�6%���U;�^�h��"�9��+w�C	ޕ�\?Dʜ��L4���֋��9����H~�c�ryIl-�G"P~���+W�Y�>��{�B�� ��M��$��w����e�a�����;����i��.�����C�hX���J�`�ڱ��a�D��]�C��yD��I�x��z�l�=q��b�%<�B��U�2�2Hk}�ƌ�Ns�ۓ�&o���R1���*#YW�ԗ��C"B|5�Rˋ��,��[�KT��ɣ�V9I�$._i�:�+661-�B�E�Q�OJ*C�ԋ^�����)5L&,���A@�v�-֭�0��]i���"��'��N�s����cC���d
bx|t�ͼ-��D�s�{c�X �KR������pM��,���}�QqQ�ޒ U�&9{\�Z�lˢ��א�����Uc��$|��[��l�ݻ*�kƴ�h�0z�_	F+8�e��S���}~w���g��s=��y�����n�/`��f�M����"^0��{RA&h_A���P<R�x��Ǐٟu�����R�d��j�<���{��d����d����2��aH��"s[Aӿ�욚�D��$;{A�����O��ۓ���VA�Lᚅ"�\]�)�e5�2B.��Uu���3=3�(�4|��#*�d�nD���Z��d�'��P��}Ҟ؎'ݸ���*�QM�<8=Ł��7�8�p��\�G����ѽ�������,)��_S=�r��q�xZ�c4����5�3,�BHO��pԕ����x�> Xi�1�1�+t��FZ^�(,�`'I�Y�͞�,�� /���C2B�t��*R}�˯�t�q��`�4�jծM�� c7�<�b[I����+?���R����5 9$h�FkX81�0!�I��1"�Y�.!`�[�.�[>��IB������ֿ�&@���+oszWb�&u2p��߾$^���^.�;�7�:��I�+�$�
%�Q_:�_3�Ӏ����CV�9�确�4%8���G�g��r���dԩJ�n7���w��\����5/e��!#��wf�ć����%b}� GAV Y�-(jN7sϛ(Q�brWJ��6S=�6Ā����V�ļ��k�]��7p���{R�"�վĠ�y�΁�G=\�>��>$H���T�1�*��jG�h�T�8��ND;,�_0������L(T}����!!ŗAY���@|�Y:ߛ_scꦹ"���������F����U��\ȍ-�N7��q@�
T==M�u/杞Pj����	�������R��(��^)�БG�"a��P��Y�d�W��n�~%�����q:S��=��ΐU��5�rS�Lɂ;�y]������QRP*u���s���Y�:����oA�z(e��F��'�����]�em�v�G9F�-q5����1�D��y[Н� H2v`��VI\��O��]T�N"	bf'� ��w7��N�.� �<8������ �G[ 0��������$�g��i��������քg^�l�ڠ��B������������9�#�h~�����J-'�!b»�[7�dn��5���c����^�F��Hے[N��v^!�������f�����?��#�qhҨ��}yD�D�7TX��*T�����c{��g��߽��"Wq��P���j�Ej�Z8V6�*�3[2Qgal]}�t�œ�:�eG�W�z*�S���q�l������U��l��o\�w�}�i���K���`
�Ƨ����:�Yf"30�ʪ�֬�!?���C->��w1f�s�����W4V�eJ��Ғ#��y�FY=�_/QB���VGО2vc��T��~�=l}&��%�V��IiEm/�$��{��֣��l��	�AxxW ����X�*��5���w��2�qι�`5d󣆫Y�U�R��UpM3�?�ͯG{x�gg�xI�pǯ.ux����SI��Z#�DTq�*}^�
���Q�̄��^�]���\��JM[���<���+j�ѵ�F��'�.�w/���-��3� ].1��S����i��������=�)���|k���Jx�6Y/ �E(���}�a��܆�
��=�V�au��2i�s[���ĉ����X[׸�X^�9���K�<����9���$� ,j���ܪ��o��-*�쵋9�������HB�x��&�M+e�Qrx�g��4� >Os�0�&�c��/�=�7�as�[	���������^�q�D?�n�3�32ʑ���En��dl�ז{�ub��s+����LX
�B�Q]������~�t��O5�s�+�1FH�B������.=vJҹժ8i�`Z&yS��u���Zǭ��<Ɋ�fƲ��[	؜�N@w��u T��X~����n�˨ �T�~
X�r�d�DO?�!�%� ���H���AĖuhվ������6�!�kAb��V�7ny��������'�٬��\���⠭�3��#O�љ�[T,��aRRܗ р��`�,����Y�o|`,�5��u#�E�v��g���#%�3�'�ߓε5�LF�HX.��U��ϋp�L�\А�� dV�������V��ԣ[v�U_rV�w�"9՛.丅��Pb��멂|6{��=(��Yll�۝�$X����,��ϐn)����0��w�BU�D3d����q]Y�x�(1���XEP���%i>R/�H��ZP;͙�8{�v�R����DMcm��Yi���Qm�Ҟ��tYB�zx�`7o��jU[|��pN��wO���C�� 2���+���}X��f����s�ad�*��^�P�%��V�+ew����z���TӉ�y��A�bKlS4ѐ 4�����*�0)�-��?��5���(^�
O+�kP(@R��駪#i:UN���.`��W<�z���ZX#�}�?2ƚ��K�rl���=�EG6���uJ���.G�o��F9c[n�ÖT��-?���������Q-�j��G����B�"(S�_$<�i�X��v��#u������0oy�
��v�\�)^3sm�R�AE��w3�6À����8+�Z噽�j�0����	�ʦU�0N�Ձ��ds�����j����qMhY\U`O��?�J�qVAY�K2���p���,#7���}�yc�J�Hj�2�m�~�.j�H>Nh{�E�V��b����_;X���
z���e3����FO�g-v��$O,�jQ�a��r���p2$c,#���Ʀ��p�y�W���i��(���[Ϝ�p�j�slk�k5�\~;���p�c~�i{s���|�apL9��9�C�nX8	L�btd��*ә�C'��VoL��7��JA|\�X�iKJ�+Y u�b���^7���)�Av��N��J{+ɼ����E�Ԙ1נxҟ&���oZ�6�ڒIH�y�??	��^�0�=Y��x�\��,���9@
N��l�c��%P�ʼĴ���b��7t�L&a�#�t@[�Z�����PAh�a� ��}���<�q� ���e��?@4ϛ��r*�0����O��� ���Ș�WU���Dvy�C��Ty�
�(���+���b���V얀W�� �I�u�t��W�7�6�\g-U��C7���F*���+�!n���-��3yH��m�M��u�^�@f��~��Me��b�Ri�o�<N�˒(�9��^�s�mc[�1�ӓI�������5���Ɉ��>�p��E�0
��)� h���A�N�إhB蠰N׋&:��	���7�cՓ|��
<��(�1Ő�ќҏ�1as2"��@1Q_��(��	*�GM����1=�U�죳�fԱ�`��̵ݶo�j�����t	� �s���f�-']�^� �!��
�
?��?���+���HoA�]�Oq�w� ��I�5��V����\�$�6ew����kU���H-Y�d����\��h������mC�Q��QrG0[^cO�o.3!E����.M#%|��'S���-}��Z�n��\4;[�H�m�\_-:��l�^�v B0FU�*�P��1p$�Ww+0Fv@'$$��Gc	�C������A�`4��U6�w ��NH�����W��%��C�2���Q��2w��$-^�Ok�<�Kts�}��*���W�������~br��F��MW��J[���ۦ�m�kG�D�a��UI~z
��&oé'/�(��� U�d	�e�*��O�����,�h2��u�N��M�,8ZZ8�=�:��ˌb����N�P�B��Ҏ�����BQ!rq�����I{­���L� ~.{X���Rۑ��@�%Mb��:kJ!�?ns6��񓁔�Y�N.�^�w��"IXk�P�Z�6oω�K��蓉���n~�N'Zx��4�`�OS5���Đ�8�
����0H��g�-�u��Ƅ�S$�om7'tY�S#U�t��[~E$}�]+̾>�.�+�/��E{"�m*��pUb�����~��c�=y�;��-!-d�v�#��㪽%��	�-1x�OHc��ꒌ�&Ĵ�����}�]l3����B,��=�飇e�q��q"L5պ����­RT^%��g
b�=�,���f)�M�]4�<®ٓ����ݽ?�@��K��aQȡo5Ҷ<�^�����~��#��~/��C����J)��+i�p�3N���Qe|x���.�v@i�5�u­ւb-��,����T�B�vO��%�֕�|�;Q	��}0�.&���E��XW.5\6	0�f����/�✎zi��ob˺�^�c;�ѡK��S/ޅ�*���A�ߑ~��B���� ;��b�Ts�-v�Z�D~к.|�`�4�
kb��5�Ѽ4,c�<�-�r�%�������:~�C���ζ� ��qe{ƒϺ�s���~�U���qN�	��W@N����|�<�"��3*�&�y����4������F�<\�*��W�����Ivd4J.�T���@�+�����l�+��_77�$?�uA��s0�� P��~��)s�E��P�xn�
�;�S+ܰ�a-�T��=��8�ԦZڸ�jTb����(�M�0�U��_h��Z��:	���,X�j���A��=�vUT���p@L����_e��M��s?��<��i��H��C��|�z��t�5}}4��SQ.��$��ĴKUS����FބG/�f���x0#$ԇ���?{�b��U���@#u�Ҹ_�l]�D>=��(;��-,Wݤ�=!�P[����i��|��9���r�z�%
�%�伷�o
���y0m�t�������n��x15��/x�����~�᰹0���{{"���j689�T� �҉;���ʷJ]j�����4ioh��r)����l�E��x���6~9GSJY	E��܉��0:��Ko�� N��Io��c�N�d�L���m��@a�����{(�j �:6���}'wK���Det<F�v�+F�<LD\H�d���XkϠ�`r�R�٢]4��[��X�6q}�zU�'�{����wvC9_���;���
y��P���*>
g�����wT�4�f��+&�NK�&.s�J\���$U��=,J
�)(�q6�W21нK�Ծ,yT;���ˮ,����R��}I��X;��M�ވ��1� ��m;;ǌ�Р����:�yM��c�����m�MI?�M��Qݎ`���%�7Av�����bO��ۻr������[`ݠ�*�)�y���M9��$��B�YP������
��/3�O��J"��Ũ���I@��%���o)�#��!h�!a��:[���]^3fD��9� �F�_��r�_C��Mޣse��5�F�'f�7˧ �2�u���c��Pl�
%/]ks�+*��nb�H���9�p�uُg��n"U&Ru�^�T�l�7ks��߲�� dΆ�F���nj��DC�X��jXY�����:�v��K�=O&��� .�cz�J��0�K���Zp7�O!�S��q����ؙ?�ڕ<����)� ���b��vv��/IA� !�@c���)������fߪ ����	la�Ll��c��/��tH�,�$��Ok��y�i���K�2_�����fG���:H\\�R��Ps6�;0���H�i�������ЗC���{<���\yܸ���+��2·x��S�V�F�l�+w��'��Tkq�|B��O8�	ɂf=5��/qx�I���24)CT��̖H�?@���_�'��3-n�С�_m�SUuM7������V�a�r��,>�m9�E⽬�.�G�>�"a;AgQxe闥��H� �2����hw$Ȝ���s����v{S_PQc�>?�a�������+�}����H{��1QXd(i���4�[��|�cꓕ��L�6���/Te�Ջ��W�귊��s>O�W.�(��T8�'(}gN�,T<ʇbVI�4�]�C��yK����[=CmhǺ\�R�i���:��>R1 �Z�4��m�j��.����{�Y���lbf8���0�*H�F�uD=�,%�&����~��sN�eM.��𗴥]�L��ڞ<q	�2	C�u�:s�9a���xV��ETۤȘ��PK(&�.��|u�AP��~��iv�`�Q:����0ɋJ����F�8�G�Ơ���tVv��`��C2ְY�Q��}A̩�՛.r����9q�`�m.*..���wN��M�Ӱ	��mH�g ��އ�u�w��
P��` %��斠@]z��v;�C�?`r.逆*���-�-/� <��ѥ%wbT���py��*2�F�rϼ]k���Ё!zu��|&���W��cҧ�7;�6#�}75T�I��s��T��k�NE"��!���P���S[�̀\�ȳ��~eL��-�k�J]k�eh�;�?�ԋ�G��(O�l9�R�`�b	�{��ʘ��+�.�Cl�H���4o��u�(��.T��>�]��\p\�ٻS{�t���#h��Rf����V]��ue���Q���i '>!�����ru�o�Wj�f�U�ߦ�m�*AVtZ��d��%�f�s����{P��d�5
���?�MJ\�t��|\��G-�����<8�G��Xq�߄ k�6qٸ.z+�m�[ҭ7h��qJ��V�����٠)�(���m2�q����kr+!�qSN����ܐ�$E�4���(YVry��yP2�JӁ��X¿���۲2�O��Q�/�]ң���GK�<���hAn��R���<�J�8�M}f]�ہMj����y�"��P*��Ј̿kz���0 IOl�ɢGj���ʻ��n��K�Ns��|ߕ�6�e�k:ibt�H��9/1��徰��:����@Id��5o�t{����O�H&��@��p15�s���R	Ϭu:���m�qsÝ�<Wϊ��A����X}�9aQdw�㶪�������U�M��A�bxV�@�YO^[����R�v �������:r���K�)Ci����g3>ٛ˨���Kä�o�Ԓ22��9?����2�BL,B��T.
�7���[��mj�=�Ơޕ��['M��	ak���9�^�=�H����l�։'�0���YE�k��������ٛM��eB#���$5�����Kǔ�ء��2�������̚be�҈ߩ%c��g���=`���N1�,��-�f�McSUG6�C��d�F�'l1�0��[���rЖ��/�
�c'�_!��ݘ�`U�B@쑣�%Ѿo�lr���-�Q�,����~���P�8�w�x;�4��f�E��(ƙɑ|7�ux�@��i���
tK"�� �ٯ����/I-�wfp�)��8��9��x����D����z��<�s��{��Y���l��c���ؾ�M�M>U�)��U)�+R�d��(a
-Mv��)�����Sz��"Hb��g����.�S4����s���+>篐� �cGlA:����3o�'w�lV�������6� *+�61V����j���QV��3}I�*=�ۇ���tb$S�ͨ�'��V�XIi��~=k�΍i�#��wE����q��4��$E�g�E�Vp�6S \�j������n1&J�Ǐ��	�m��(L�7��]�^�$�zï��f��LĸA��$t&ј�'�̨�YQi�("m���3�k�I�����o��s|קi�&����d����&��V�7��䣭5٥�BaG�/�U�憿��萛g��\�QE�,Ն��Q3���\ԗ�>�����Wu4�e:�"Bb��ELR9���Q�L4�u��
q��пk�+(�k���gMa��.F!�+Ykw���4�ݱ�Av���*2��xx�w�$&��4K�H|yV����q�;�D�mdm"�t	���xMZ���0���,���[�6L�]�ǌ����P�n�=/�F� ���IirS�<��M~4�;#V�p|�������v>LWI��,��d8xAW��T��]z����L�g�Y�ͦ���4';�.�P�s7�ou�ଲc�B�~��}������78g���8��Nl�+�~sB���		�7 �!�8�����W+�ȑ�B�]12Q�8Vp�=���q+?7S�|�dBE<1��/ac��RsD_[�����$N>��g�Bgs���4�q����*��Z����6U���	d�#��L�X�G���6>4��}�O��&�ݷ`6'�7F��9Fw�@H���)%Kv=?��hq��sނ�aYD��8�I5�X��>
zz�,$l�Rb��0�.��ޯ^���)T��;
B�1�����
V{9-�z�\T�� y�ţ�#�_����n]����m?�ֿ@.�c�j�prI�72�>���WuQ+1OH�V�U>�ز��,��2ѳ�fL*y��sY�W)��A;��KSE�;X��ba�����T{�������gɉ|��ѷ��Rͼ���b͋;M���6�E�7L,�i�i�g[g9:
��}s/�O��A�WՀn��1yc,�L��r� ��[��꺻���1Q��"���W�uv&���y23h]��9�T��"��6���s��z�\�[�{y�}�K.���7��(,�%z�����	'su�I30ߌ��`���Q��D}6I.�߀36�_���oͫ�4�{��>�A��{��Ƌɹ�~��)�pJ!����D�/�re�[~����p�W��Ox*�����������`p7Ɏ�h)0GnY���pP��8� ��g�(��*śb���nd������1�U�������ٛ<�B �Y0k�;�X'
�-�m�k���ػ�^��
��,	"��a����ɘ~��M���Z�C'un�o�m	O�������,M�u���}��+���{�����\��E�KJ�bu��m%���/�p�q�iϓ��7|�(dy�7$y��\�Cf;l���H
wt�6rO@gS�/aG���dJ����ٱ~����x��{����G��I9��j򛘣�=��2-9ny����{�vЇ;��D�K�u��:��g�{!��(��m��#�מDg:�"Ś�C�f�<ȟ�X�"��dB���65���p�>Y�Ѣ�Kyɀ(f0y����ѿ��8�)�6=��i䨀�Gt@t.OȮ��֬��V9�ȴ_C^���h����nq�i��_.eU�(�ʢ�!�*l����\�z�vgt1�X]�W}5�ޠY����;�ݑ�B����Zm;;��M<�,7�[X����%h�܆zHd=Z�	�Vu�;���
f^��~gU�����Ɍ>�W��^l�[�����7��n�/+��&?v9��d��+辇D{��`��(�%�L�x�5�-N�����m��V�������Eh��SyqaQx���T�gHO7������Z�?1�H�$� ��:�65�?��#J:4�q�a�W$�K�����E���o��A��V?]��X׬�t����-���$X�u�,݅F܀���;]���x� ��r6�Z�R��?{���[�]�D4�f�$�_��l�B�64���᮲4���
�Å���]cJ�As�N����#�-W`k��Ӈ���H?�iF�����%�.�H�����>����>����1̓��r۶xTM���6Ё��&Ц5�h�[S�2q�m������4)�=0�8n.�i��D�%�����eGd:������5=ë�V�5���,�f����0IVv(� y\�NJ(x��q�v�G0�	�<'�����q���5+�|�>k�@���S�����h��?�:�X�_�+�nV֬.��^>�A+��P��	Vq���j$Lb�՜*�q�$�
X�X��1��/Z�b��BA�K�����fn|�ʥ��^h�D�ڹNagŝ�����?��k��s�p�Ja�tS��/3.pHV'�K5��^�Z����l����������pR�I^}$Wx+�|��Ϻ�bMr���Y��a���c�m�����~-��:�G߰�p���e�w���"��pKP�������¥��q¦u�M!q���|����II���5�iJ���d��'-e+/��y�孓g�!	Yu&����I-�ԑ];��4~�A{KȚ!#M�Q"l��`�=%����7õn�̒�F��f0�U�:�p�VK���1n����7P���;6�DV�c����LF�r�#�C�cl���j]~E��wn����i�I���x��eP��5�m�TL�w��U���B,������9|������eި�a%�QA��Aړlؾ[
��V�v4����]["�6wR�j�uk>��LUdΜ]U�j:��4z)��d��>͖�����VQ�;f'����n:�T�^3��o��S��pk�X�NE�b_,�Q�2�j`���$� �ڀ�<��K�tG�ԇ;L��p��V�W/����RVI4�ؔ *���)o�-q������H�{N[W��A}�>x��C4�ʆ����>@g��up�l�P������f�����˽�%@��! �R�Q�^&�Z`�ה�b>=0�y
Š��z#c�V�Ċ�&M��`��H%7�,�[o�xGxa�YCZ����9�_td�n�����e+qӋ�6M[��+(��6:�u�N�a~�_	L�ϖ�'݀���cTw�O�'�Y����-#ڏI��T��u@KtW��� �d�+��(��/��%yz�zm�HU�5t�WN �Ӓe�3�>vGH`�ɍ�f�V�ņp�?~X�؆�h��#��e״��E���q���k�؃GD��&����h�?��"������<���������"��}N��p7��� �ߠs�%刴���R��U�B��%�{�+�Р�����r|O�<�F�\�Z��ʱ����{��2�<���I����+&۫�WzU���t����al=M��ʌ�{6�E���Yjl�[��H�>n�k2�E'4�k��Gq��~ջ��J[ַ��g6���8Ѻ|]��Lm��O�`�̐�����]���t�z3b�'�g?~\�0^��^,Ნ��o�	��C�h*̼��-���|�R��1x�ř���\��8J7NY��%�LI�-�0G:ך��B�lR�'�@�����F4L����)�q�5�+z�%�O�X��\�#�~S(eHP���xN�R��Ǡ��8�kg�G)[zBug���}�_^���{����0�[���+;��9�@�frT�\��iJ#��g�����a��+͌`FZ���{�Qu�����e����@�2'�׉�0\�@,�x-�H���AF.�� "��T饭�5���H͚<Ta�m-`V��xʫ�XQ����d����d���%�����y�(Y�zx������$��=��� e���1Bh�\�����?��╼�^Q���EKu��A.=�����%Qs�D��A/���4k[�����j]�A2N���LM{y�I;R����Q@^�<*��|��ok<Q�f���]��X��5����x��Ϊ���A�K_�� �_b��K�$A�혊����d����gN~�q��V��\������H�w40r�@1�j���TBZ���tk�j�ܘ�����R%�:	 WKG5�V��������l�x���O��������r�l��dһ++���[�X2 㝲C}B��i�I#x*nnK������?�k|*"/��s)d�t�p����ӳ$׹X�i���h��u���4��^�ʟC��A5hU1dg�X�A��hr�cZ��t�?߁�[j|z3P�4���:�x37Z�^zt[�'�
�5���>'�X�{C�'eMl�R�M�����c�z��+��ʝ`���\�@���j����.�x$�D	�AF��t�ަm�D��%R�,�]���.:�#ζ�{hl��:�LI	\�2.=�,Ւu{c	n��a���Is��-�'?s��m\+���쐣n�h����vaj���֪~{B�q<������Ɣ�����c ��+o���6xq�	3�J��%�^6U��N��uҕn��>��maW�ˎ�a��̿A���M�����F�����u��̳�S?gD<_�N:'��D�)��1煜V������5�j��	�S�g¹���&o-�h�� @��N��E�R�9��q��0�\ג>�w�����)�����>���Kt�U�%�ѧEikSs�Y����V;���Ц3�����#{��������a<�'Ҵ�Q���yXxAC9��	��c%R��@Q��{=����h�N�����E�^��	X���s��Ā^�Fm6��3t���W./���LTq�X)���$dJ�{��6@��ֶ�4id楤�������\j��D?(��_%5B��,U3��h��!q�O�d����J���EHh5�(�o�>ьj�A%�SS��r��')�" ���~��j�)�\¡z�`�>)��AE(^N���貧E��wخ[ˇSf
��5['�n`��ߒ�%��Y� &�w�&��3ɍ�<�k�)�7���ʎ)]!��7Zu@,zZ7�ܝ�'��P�ʀ=�O�):�Z|�q���?F���D�Y�E�z���dn�{P�ܬ�3�xL6T�ֆ�}��[��۳��v۽2^a��>8dE�Qv)��߳w��3��ge�[����?2X��ɂ���J�؎��W���j�w�j��2�GYPy�D��Q-����b��~z�����g9ڬ,���T�^�&����3�#����H�w���r��ɱ�Ჺ��z��:><7�83�CȈs}�R�q��,1/�)jW�V8I2��/���Ѡ�Ϝ���L�"yb">��!��Dd�]�{�d9�X�u!d%��Wdl�7qN-�Ŗϛ�����0	�'��(�N��fE�_L����Qj���8>��8��I2���7Ay�[���k��T6 �oΏD��ȃ>�O��~:�m<�n�}���,C����vLo��� vj�h`�6B�yƮ���Vd,pSN����W%��$����u�ؽ���b�G��*����M��5GV[���7Bp��˺��`��~���x)bJ�9[��Y��OQc?q���Ҍ���6��6����9mS��<�4��@BG����~6`8�T
2/g ~׸�F�œ�U{�����6�@P~J�4H=a4��S(X����Lg���m\P���C�R2�c�^�&W�f&�1T�l�C]2�2���<�����ƵuL)�P�p��Ӗ�K\�F��t�)G��<�!�U07���i�Dp!��}��Ř8G�H�ŷ�������,�j_~h*�𰑬��#�������s�G���9���b�C'��`N`<�Y8/��@���YPަy8�l�Jв�>�)��	|	(i��FT4�D��|o�N]O��!۠���ԕܗ P��-Y��Xx&��&��գ�`�@_�/_cwDEGlfMw#9e�&����J����%��t��-��w��6
CɌ��C�H%�>;x&mF8��ָ��l�H	�e�uolaێ��i��w�2�ZM���/z�B�'�w&K��
S1��7�z"HZ�`�����VM�WTی���C�z �,ǣ�(�J�/�zB�0Υd�QeЛ��+�}0���2[\�	$����9�H�����j08���R_�\��Z��~����7K9j���EIz��2s�:�d?�(*0���ZF[�Dq�ր�,�����#�Lh8Gt��\��D-�p;i��η�F�;��/�k�6�v��d�L���HD���,9g��>�?e2e��5���uj��Y�iF�Єwi�E�D��8�\e/Q��}����-\��A��?��x���;�kg(���n�u����
G��,�Iƾ�^���ƺE^OXA���nYר�Pb^Y�	I�M@��AL���8�[�r�����!J��~�Љ�{�i�Z��vQsH�WwZA������h[��IO��������7�a���4sL;Y_��a�� aa���Qh�����ݍJ��M;4��E�[��X��me��NՈ\�}io*��U)�N�k��qY.���t�E�!s:�لW�kj>D�o�-�AJ�3B�#������BT઺�n��e�~).����ƢQ�x�,[��H�
�1�F��,�ȯ9[
��D�NXS=�e�C�(\�S���W���xN+t��/�-B�.=�UW�-"��@#�nmod�Ǆ!l�8��_��έ�����hr�GIZ��!%�����ne���HE��bo�U�5fm��m���s׃�*'J!�!�D��\����eyP����ة5*ȵ��>��[����ԊP����[�6��be��v�u8����/��9;��y�B��q8I�]!��
/�(�x�艒�� �����Zl��kp��H��zG"���5Nw����U�'���ќ	ø��M�)��G��x�%��׊�R��ku<¯�{�6U7bƥ�m��$�@7Q�����E-����<�Z�G�ѐ���e/��S�&P����&��.U�������>sa��Q�[�\w���?e���=ï�hq,��nK��"�%�*��@VT�]E���;�`�rub�у��0����*�j���P��$�O��'��)U�<aJv�;SZ��ۣ(w�Ri�h)>�b.�c5�@��	�d����[T����gw��JmH}�%�h�{'A�����|��z��6"�}�������b��P��ML��v�.,h��\N�-�B9��_py�#]d~(P�����O�Y�x��c"��_�0���#0�ʚ'���y@K�8�����Ǥ��+4J�
řB�֌�����|�K�ျ�ڛ5z���!��V����WQ�F�����u�>���ޅly�0��:�������ڄ��×$j��)郴����X0���*Ї9��F�_���D;��DU��g �w���{<���"EO��g������g၎-�}�p$�Z<h������ ��>M��At	#��򘣢y,�(,�����ǐ��E.��p��S�:F��a���F٫*>�&�V���tŰ#H d��Y_�`u&�0tmO�Fa<��K���ZA<��Y���d1ܗs��a5�1eh�i8zؑ��%/&�N���S�/�l&/�M��G��Ȝ���+g���n��z�SŞ/z��r�F�T]��O��D�~fٟ�g��Qe��u�k��"k"��sx�T5nZWY��BQ��S����gJ�켫zC�~Mʑ�P�:���Ws�q��`l���2��A�J`�3��z!�j�h��)5�΄��~�ʮ���(��q%#��"[Sd+�=�-h7AEy���/㏙��_I�WU&J���-�Ry�F�4rc�� @A46�9�fM:TS8 ��s��;�%�8���]���V��}1���7e`As&���YZ���4-#�;�i�j�5n7��p|��Ma��b��:��2�;���i�FH��(�^xg=��Ş��CȷyG�^�']&%x����y���b �7��ٔ�r���m�����њ�P����p��+F�8V��v�&�̭��Te�[a���PQ"hY8W7y���}W�`�m���M犉�UH�u"Nzƿ��z�QC^&�hݱ�H�9> K]����kف�v�oЦ�0�Bj�C�:@��/�\.��`�AL��3Ș�Ҝ!n�c�0E�����(|
�v�Bs��2�*Nu��
�t�� @�v�)��P沎���i���$c+=�b�VuԎ�z*Y�����j"4����Ы���A�$ �6��}�7u�>T���?4m�5t��T�Ҽ*�S*����"t�C1��<0��"}Ҫ�L�p�P��Ż�g�����z�Ɔ�Bj In#��ӓ%�S"�?g%��ث���#�a�r�G��ܨe��.[u�S�}�ՀMSUk��Mp�t�xS,MD�m�*`�鐡�����2�`�W�E�|��:�F���@���Xc0��A�u}���B�1��������� ������j!��ՐڵY�6j"��)2�K q�ǫ�[�Bm���1�NF� �"-���ܖ ݬf%�c�FסC�@i��A�K�lԖ���� !�+�''�䌰�	�\�T$��6c��5+���zr�F�3�E;@�4�T�Z5 ��Q�����B�Ɔ����[v�w��6՟u�WH��Hi�AtGZ�$��_H.dm��}������uג�g�ˢP"k����/Cz�G�*):�<[��Q��'S�M�
�y��Dl�i �Bj���3�ndvژ��_*�,�b��p��k��5�t��
�伫��R_9�)6��c�� [ʞ����υ؄�We1�/���e(���m����;�Vg���?ω��,^g�u()�'6pm�b��r&���|���>��Qυ�k�˭I�1��^��j҂�p�h[|4a�*@��+�L�'|5��1��E�d�ڜ���z}>���_&�V���;	��k�T��ɉ���� ��]C(�g\P9�$�J�awԊ���n��Ÿ 0���9{¾0b�`�cO
����ܡ �7J��Il���<����;M�q{k����+�A]Ӝ�_��_�#���"��@𐅈	�/i�����Ż~�Y�g^$q�z�Ӝ	��DC��msu��KJ+��\��F/�y����]��&�r�*����`2�M�6�f��ba��GM���a��Yk���(��~hx���=%~��S�=�Ԉ5�� Z�`Rhi!-'� ����厍�oqͱ�M�sf��J� @��}���D�R�Q�M�5���5Ϛ�on��{̍@�VTՠ�wD�Ao�`k�*���xYJd*'�-Xq��ŋ�W�d�IJ�r�䑨����أW$夛6��oxA��;�3�ʂ� d����x��`\�|��ü��(���A�"z��)qtTg®�f���"e ��S6͖ �7���f�A�杲����J�͎r?��&^gܙ�Q���d$��?׹@V
gT�/�� X�9Bc������[7aM�hq%d�(���Dɑ ������pw��PZ'D ���R=��[������¹�ۆ�y��?��.?Vo�M�<gD�8pG !�5F�\Y'F�ly�~OV�:x�j�cl�Z	ͤ<;w&x�Cj���p��L!��w��,�l$W!?pQ�`zp���>��+ ���`�7<=O/���"6HY��)�+%M�7�f/9�k󔙕��T���H'� ���|t=X("])*8%���}�Sc3�b����{:}J����!U8�~���&R? ��QR�g��ZR7�d��&���K���.�)�7��R�Q⃅��.!�3?_�R!�U(f�+������}peSqU���@@�|�4*B����?�"D���]B�:�F�#���cv��Kc� �tSEx�|ml��%O�^�
���(.{�p�q��9����a���R�[�D�Mmb�mg��Ժ^%Ok �IL��Lj�Z���@�nrO�>�-����|���v�y�_�.q�d^F�1�⵷:8y|���� �x��WVѬ�t�'��9N\��O��L�g������\��h/)��WIc۔L҆�:��U�cx.L0A̈́H���Y,�� f�*l���^�m;2/�M[��D*<?eFbٵ�?��W�q�Gw ���P�@�)S�6��AU����|����mZ��E���R�I�[�"�y�fk��ѻ��Y�ɾ�A=C��x�]�w�Ca�g����,F#�#�ka��g�����1���䩫Y��"
��'E��[3y<��GbV�9�$ooGعY7U�~p�vP�/��n�10�H�ܳ�(t�i-1��n�����>�eJ����%Դ�!9���t�u7Dò�!Y50?Y!}!Ú������f����n���$Șe � ��h?۸�0�p�Ň�[4/������S��z$��7�N�V�?\?(bk<�v1�P��Aǃ���9W�� �W� ,�1�W%ɠ؃X7�%ڵ����[�\	*�φ^��D���^�!��̾�_�1���Ѫ���4�Z�B��x+�;�/�rW6�J���T����x�!���z�CͲ�� w�*8��O9�9�g��v�e���WU� s9��P0���$⚪��<��u�V$	 ����FGh��@ٷ'�O��; �z��FM'X".$�-t�������S���^��-y�2쭹�$J�V�����Q����{ˋ�Qp~��������G�\�6�GHt�6��X2�ڎ�+)�G�v�] �4FSU`�	� G���_
�1%��V����X7 '���6�u���5�tF�^"=sg�)O�|E�&�(�'���FB��n1�� l��L�c�B���	_W*S8g���"W��"}),C�F�@��|w�,�o4�
�r����)�$~!u��Ra%O?�ϛ�f�h��c��Z�$Ȁ�Q�Ӽ|�����O5x���>��Ү���)t� ��%`kq���4�.��V8Dq�`[#Q�[;ў����Ր�:(]���(��`��s;"�o$*���8�cP�W�
����A�k���	y�$�1��^%����������c�f��p�Ꮰ�"�PuP�v��6	����!9;��G$��I� Pyr�6U�¨e�ni�S���%=�M��R$c�ٹ�-�����=����J=w�:��R��\�+>���#-��m3|r��ǚ��No��Q�,� 'a~��/��$�����=Yg�&zs�r8�:B�0��h��R��S�t�[��d	���)�EtU� �0;l6c�J�p�͡Ar�{�hj�ڌ�l]74i��F��6ɏ{H�{	�;HK��4�[�)W��w����O���� ��5�sfg-��u�rϟE�e�"53kr@|���v�p�]<A����0���*�y)l�(#j��k��;3�& I{ZSg�p���ʅ%!�S��=g�Ґ'
o��A̫�I���UP�V #:*�'o=m�z�?��Pݰ0���q�u"vps��&m���NC��O�� gp-����)��1�Ѥ}B�r�j�7���1���2J:Q����͟��O9���7����8(e���?!~/]�. �YO��s�������g�4�j�����U�&����8˯��(v�ɑ.��E+��~��8gF�O�sA$f�߁kG��7B-=6�^��#B��p�~|�T#=�M��}y���{j��`�JKM���o�z�~���,�R�P��K�+{I "Y|,Ǆ<��{Q)I�DCC�Z<�l��s:w�M�q���sF9ֱƖN����F!@UҺ?�D�}��;r-�
���Ξ�4�{����7��6[�j��9��:�l�K�����ze��W7%�T��(��9����1�2`�1D�FH.tn8jb��#<��dI	{~� �@�]ly�]L����Ct�Zf�"EYե¯�㎭c��rR�tp���՛NC�/2��E��W�������Q��ғ�w�޺�}
Ka.XqI��
9m�N?C�u���&��Ѭ��� �a+y~�a�8�%�U�_!���/3:IC`7���i�I
#�O�۫BI��cJ��G��<RL��0����k[��������:�A+ի�+\^�un����e�!�_���y�̂,�	*�Q�In�R /2b���WYe���w���QV���7�<Q��9r���b�&�(��WO�~U'Md�S�C�T��e�l���	�.w����iH v�آ�R�Y���F��7 �㩃�&q��c�D���Aa=�!�8%9I���˟��t���j�mV�5/\�Cd B 1M�l��4��$�sb���۾��� �qu�z����`�"L؜�)|ʨS]�WM�=�n=�?�L��S�(��*Wg�����������o�����حN�b��?�d��
����Ȗ;�p�rZ���N�q26\���{�|������{ܶ�I	�HR\aW�����f᷌/P�[��p=�QhH��i8Aq������y8�
~��C�TX�gQ�����v�6ö�����d[�w�����_jV�\�݂�%�I�L��Jq���-���|K�!�Kܺ���l��ڧ�e֓E�H���G��,���b�B�栨�u��������������C�`q67�w�L�
�&s0ʭsK�������q�M����y�<f������QGj���]@	m�=2/���	�Rfjkk�>�b��ʩٞ?�%������[��`�K����~���+����2ۤI�t��\�Гm޼،40N��=�oj�؊z�|��⌍V�M�&C�
tK����t��ځ
ų�)�xSXGA������Q�J[��I�!n��ɤ�`")jE���YI���\����U)�4 ^7;��W}�����TX������#�%#����k%V�c�-�]y�K2GN��=bv��1[Tϲ�/j��B�`�jQ
�%+�Hb�����4�E)�N�8�H���t��8�+=�柙ƹ���sH�MdI��^�k��������cVb[�����56�z����
�+�L#-@���\c��f'�5f��� 0r�/�eF�O��*��9qA���
s��F=���m�nA�IɽvP�O<��y[crF���,y�v��j.6_:R�i�Q��͛+@H|&�䴩��<Yȿ��6���'��`�l:��3�x�ڪ�NL��&h�4[.� �\D�����
�U]���?���3�+z�w7������wj!�[���L�ϼB�JF��u�%r����vk�w�w<H�R7��(�ASy�yԁ܊^��ƀ���ȋ"��u%�L��L��&V�����Z�◧f*��@Ȯ���n6{�p|�"��Y���	.䠭�J�Ρ�]����Rzl2�!��i�dl	|f�]�ͅ ���O��UY!� �t ��Z-O�]�s�6��'�s��~9����U'��xSm�IB�Q���Q!�Q��ן)�a��1L(�ܘ�}Q�U��铄*V��?`������I�e���Tާ���Uo1~1Eq��F~F�n���G�j��ùJ��:�E<Qu����p�`2#����4�p��'g�3�6��v�D�*��hB�U���0����QU�:��㌊s��#�����;@Һ�Ǩ�/��Uȡ��;2���0�҇� ���ێ��N�ƭ����R�K�2+-�	J�6G�(���2%�y�q�G�wݍ� tt�Rs᷷"�.}�Yq�|���e�����k��c���"��F���@�-"eΣ�Q���y2�q-�Ye"����DD������h_�J`���4��yv6j�Y-L҃��*�9[d�ˏ(SP4���v�n��wc7SwLh	ې.k�������QR�#5��D_�*�wP_j����~���r��y�{�������9�
�ֳ�����a/��,eQF�#gP�V�\�ˁ��������w��@p�4���Ymr���L�h~�X엄ǥЅ��k��@k�9�KBG�=<'��O���a�� 46��'w��`*s�Jk�%T@��&A���7d{����O<퓕�U����ڹ�q]�[�h�g+k�ss�y���`V#�R���TO�Z�T��A:o?+@����Í�|�bK��l����E�|`N��lୠs!(�����od 6Y�C��//>s���)���I.f�m*i��X�,��d�6�������l��!�'�6�wp!Z��"�%c8�'���r�!5\�LS�p�>�n*}�fy��4���t��o�ƒ��F �M#>��ޖ���k�"�d�m�x���Z'a����u�P�I�B34G���$�|{�ISM
#�o�-%��µP��|@�ɏ3m��w�\v7[��m .i?6�	�ml�*��4�/KL��r��������{���W6��ߞ�]�RT\v�����^�.^bŞJ�%��V�%� ҖS�w� ��'��	�㻭�h�n�f���|���0/]<��<`]�1�B$@�^�.G�p=�(E�B��zi%������c��i� W�
;�6�U���vѩ��3ڕ-����uo�OT7�Əo?��WŞ&���Ȇ�d���� ��j_`�r�t+F�O����#�}tHAV�(�C�^s=��<�`c�d����S5������6�)�ǃЮ�W'�P��1Q%0��`�ޤ��-ܻ�3$��߫����%O2����ޙ��_� sçLa�6H�ccn�
�nIO�V�yg���t	,�i�C��"�+�2�3�-9R���ţx��}!b���S��	�ՀO��9�QkB�Gq�v������QF�Q�����~
m�g�X��ة����������;��.qw�5�I3U`��d�9�$����2�?���=I��e��A�.l7'ɦA}w*ҭ0Ob��_w�{��g��BN��P���Ԙ�"��Bj[|p�>�Fq8*���#B��Zz�����R��z�?d��=<'���O7�s8���a/X��kُ4�7Lτ̛XZ'����/����n�xvO�Z	�@�wI���3�8�q�|*y�9��xBO�#�^���{�7&�u�����|r|�����b~��/�
ay��1�K�1�^����5���x�j�:f�D����P�'�<gQ6�b���S��|ie�)b�ݓW�)��Qaj���<��=b5<AQ�|.�wA�qr�׉g���u�Z+)Z��ݨi��=�t7Ҷzo��$F+�b�7<�Z�H?2׶jL��W` �>�d��[�&�Ŕ>��n� �+��k�aD���k�A��3_eNGL6����� �}�ݷ����_����y	�X	hV���j�71o&��l����G�>g?�[[��^���� N�;��m8���������^���>�i��$\��Sa�����>�iQ��9j��.���s,�k�ob�κ�r݀�,M=��yk�X��-w���g ʭ�f�����چ��U�v�_�;)M)ry�w�t��E����b�c���I
ϫsi�=D2����Yvh�s������x!��c� ��n+��'��{Jؾ�����Q S��:�����9�l�/�w�z!�̃{�9��]o��Q�N�C������C��.ea.���WX�+z�	݇���f��)z]QE+z�+qY̶)X���������^	#��Qo��ĭ5u�?��wm�0��S����*�����Z��%�݄y)^��
�
�0 �էA Hs�yR~F�{�H�m&q�8;`+^Gv�",���а��P�e�Ο����VCqуb�E8��OꍠI]��� x!��ee:2ֽ_�%`T���H?[����++O�c4���gB������,�t�YW`ڗ��^jT��w)	��6�=ȁ�� ^e��1����LE�8��7�����Y	Gf�m�
�� �����.�V0��L'�}������F$!��m�E���\����@�]���C&W�:���}Ր���_��"��-� p���*��~���#z�,2ѩ�?��#3o��N�(�_������L�x(��VϤ�����ڍ�3$ֺ'מc3{z��Q�ׇ�[�K�钜M�h�7?7"��Å=V��6Д�JΫU�'��*�WF�q~N0������a��a/{����vJ�*a#/�P�gw�S�3�����n� ��X���%���v\�en�v�
�����6/,R����YI�AԌW��@�e	+� �=<RM���o�BW�Og���#���l����v��1�K����8�����o�Om��~��0�_=֯L1��ϟ�-���LiT����=ט6�/yG��+BR uO,�ql?	�sM�'�Z�d�]�T�=<�����5S֎ޝٽ�A�G3*�=�[<wv����F���W���y��3[ZM�������u0|�B	h�:*�)��Q��CƲ9��"żkć��sg�P����J����Om��������^���?D�bh(чz�m@�TP{��൱�?Q�gDDj��!��	��z�l��L����i��3P�KW���}v"�6̍3	;�u`��d��"�X�qjzk�$�n�q!���2�,q�7|gT���Έ����yY�\�5UƩ}�/����E��|�I��6� �Zo�4��ر���Tc)��T�*��6�\0����Saw
|��8���ObH	&���.����VR���,�m�qa �^�X}��DB)�%4о^05�����N���_�����y1|hm� ��,h�0���� H8�%�)���U��M�n �\�2�1d}�!�&��6�I��q
H<YmX͙
��m��� 0ATQ�R?$EAӉ��^�p#�K�p��&}�ds�\�WtX����1���M��uy��0z%=��鍤)��0ge��ͺ�ݲ5�������R�4dA�b0 �WH�0��i���޵� 8(�o	�tTKn=9��p2����}���Ǽ��#ü��V>�_3��jp�4	<�y���p��y������hZ��W ��SR;��
U�����:7v��0\����JI�r^��1*��h�����J�����)�G���L%C��S�k�2
`���?�𔧃��\�☛���na�	ߧIG��޸)�p��vh�Jj���1��G��{6��E7@������g�y��)�U��3<�ǳ�v�>�v����Oh�9���`�ǭ���(3��t>Qjp�0���C�0� ��Sa��DO�}�"5i�_��1�å��0'�ֺYs��]""�Y��)2�:<�ζ���n��9���ѮH��07E��p.\r;Nݿ����Ź��@�6l,���Cy3QL$Z'(�L��hd�sL��(Je���@)���4��BZ1x*�(�?1�Am�D|vO,h��_^Gq�{L�տ��>f �u?:	Q��I��vԓO�1��|_��A�l�5q���P˰�8��5S��3H�ċj%ͽ*�p���ŽǤE�� @����x|~13�S����h�B��n��s*B ���4*�k�[�hEXa����Z2��� �����!�L�Ϲ�����i%V�2�������P��*E�2��:n�HM7����;�]������V�,K�ȶ�ˡr	��~d"�t���B)�u/�œ7s�G3���D99ʷ���D͜ѯȩA�s��{�g��j;�'T�����U��0�%�����W��a����AQ��eFp�W�G���!}O ��ܲi�?�%Ӗ��J|��8p*$-�����W�8|@�𳲁���#�*"�����A��)��X��I<I���t$=j�ZyZ�"aT��OA��,��Z�5i�/�r���*O�-J�(Ͷ�ƶ����Y�B�9a��IF����66l�
kn�-�M�EM���K�?��`�Zr�T�n�$�$?b�i���8@H:~![.��ʫ�*]��������VA;��
��.#^S*�1b�P崘i�A�h�f[|2Ŋj2@�>�����(m1�)^j3�>��B^�X�]���ܩj� aZѯW�O�w�xt���=#�q>j�^��"�U�_c�)�#�Y����˸��L_�A^� 3�w���4X������4�9<rcբxWi����S��ƹ��f0ϑ�x���!�ϣo�_�)+m�Pv��ɼ�����g�<�/��GҤ���K��P,�Q!�G�����˪;E���+wS���i��;�[�l��^&��bpBq�	�#+�����}���Gv�_��z���i��`09往A��7����d��qe��\�
��53/�w��V�H\7���OS%c��v:��T���A�/o�!���1P'�dH���E��A��W���fU�d���z���K
[�G�:"��\嚰a��߱k��ζn��Rl��/�p̋ĪZ��@ی�(�1�E�N�0�k���'h{����������L��� V�3B�$�p�|QQ�#Nq6��7���?_�0�B'�6jS����@h������j���,�x�� W�]��ō߆8��а!)��n-�Niׯ�y��RB᩠�}����,RsҸ`�(�a��՚4�r9}n"��n,3@��W�D��-C���#��jB�yZz�1�D�T� �ڤ���#Fw���ͤ�Vш��a�� ~2���PܳT���]q���+$殅�#=�H�<ST�4�"��i�W�Pko� �u߮�~�2��H��
'���Ji�7`�I����.Kܭ:M�bXD�E�i9I�49;p�䞜�S�gf�{gu�(��3���ݚ�P�D�Ǩi6kZ�Ȥ�s�%����z�"a��ܱU^��Ǻl���ji��#9����H�$�`��.�<��X�p ��5C��!ECl�j�Oe���ݢiH`�q�����'d:uA�lq�!k
���?z�!틿2�Z�ݱS��Lhb?"-�H�?�������m�	�*w�s<�r$�������"�{��S�2r�+ �OoU����R�W��S�aͺ��;
��%�|_p셩�߉�-J9*X�O�������IZ�T\�s�Z(FU�#|vQZ�Qe��@��7��l����9W�`[I@�$!�X�֙�!SIZ�n����cG�E�E/]@��1l+ހ\5���鞉�s�怊�
����z���!��,�����J���{����8x��w�}��҂yX1U�E���iU 5�4R,�N�!�9Z�(aB&�Pb�$ޣT�6f���|F�.�*s���;M�0��U����<ҧ�9�&��S0���ځ̖1&��Rwj�Gpq�}����^qL�Ӊӑ94��i̯>�@���.5��o��^�<Vӭ'?O^̠]��W�4��b�߶([}��0.c��k��N��}��k�y �q�ܽ�87
�����A$m�3�����Nw=����ͫi0^��TU&��d\��`3wᒤ!iH�A��#�j�|lm��\�ځ��֐�b3���T�k�!�&�qh�b����,Z!�Z���k8�;԰(��uo�D{��r�A��y��PF:�m7.X�żj������/j\%���Q����x�4�%9�+�X��nF~�BJ�F��b�S,T[�țJ�*�V��4��̎`ّ�B�ĆI��5���k>O,����vQ5�>�g���6��6͆�����yk��_j����5��,���pk�L�ܜ2O�#>tCqU��㔖���3Ұ��/��]K�S�4A�~�����#R���Y��:a����7���;&F�����-�����I�0$9@�[^���Xy��i�q������9T�K��Z�@��/ԉ�١oqogJR<mU-��G���7Fj����;c�`x�@���o�SF�U��J�JbgE����1� �M�j!�}����콠�Rg���n�[x.������E�z��Pn������o2��@��m^�Ԧ��
g����qL����f`�b�$>��ҡߴ��^�XI*�� B�}h���xҰE�����(��STe��I�x�4�t�4t�����iQt~/ ��:�wSt�!91)��H�LEC빕��b���=�w>:_8[�x�Cd!@#JU§_�J׽dԘڏ&$bm�Ku��̫Oz<�M�z/�8{�}>���Zt���Y���d$�J�ޟ^P��������l��2k��̩�ޤ��. [���c[Pl_�Ʈv�[�׾���U&0rm��?�����r&��MD\�еC3dv��G��(�;�����"�|*�{{�
 �pv����C�����l'-�'X$I�Ɍ"y
���T�B:���x���Z�n0�lhW��}����4�,ze�� �͉��C��LZ�3�i�*K�Չ��o�E�i�Y9�ڏXMȼ�"��q�3�������S�Ie�{�w���oá�K-�@A�J���8Kh�j���Xs^%z,5�z\��2�~�m}*k{��Ye��aE�*G5��:�_x�(*�,����*��Ȥy�H�m%}��h=m���2G&s;�[c^թ/�8�C��ubd�,���*鿾_O3yv�7r���x�����ku����J��-|v�͟+��p�����\u@윢�L"~T��c��Q^��N���.6��(X�q�n>h��",GJ�5���՚2���}Ր�m����t�m`3-�ζN�q����Þ�@��(P�A����LΜS��L��.qJ*�jB�Wg'��_���W��'԰���Z��D��%��ߥO�$-�t��4O��m]|��׿��HY�NL�C��5��?�!K���6�G���")��bvKb"������d�"�%>�-e���6 �3���C�Q)Jcx��|��y�+$$+��?�\���'�@� L�
�X��u�e�r?�T�/����x�J�O����ޓ��c�&$�ģ�z(����̎7u��Y E��n3����U����^��/���t7�#�g�ϡi她���I�oF��c"��bf��ZT0�����B՝���������ɽg>���0�(���aY-R��s\�E H�=�C�,*�J�-=U=��~�<А��M9;?Ӄ�����$&���������h*`�:��i�Ozq��3�F���>�M�}Xj�Ah�U5�Z�r����*�
�W	�ƥV������!,S�{�xT�/0rS2x��jUSw�A?Qf�T�h	��*R{X/_�?���{��'�vͶs��`��-�XR��C����U��5'��u2�Q���v���A_��T�{�T���n&�������%2E���t�����\�N��7;PF���.����;�����-e��'�uK��-��0�T�f%���y������lA��:2��Ǻ~j��޸J�m�^!����t&zɋ^@k��4�-�Ӻ�2�^(��pe�F�N���M�bO+_��?X�5[]�݀���5��D]&�N�`���!�D7
�;���6�a5��)��@\��Z�	�RsӖ�=�^�9�1�St"i���pu3u���#i���o`a���@���l�.6Ҏ�{ ��S�.,]\��9���T���`�3Q@:E��}�� �ɣn����,P�X�+��jb]��Ȇ�0�B��}��H��o�W5@�PN�^g�e����<Lq`���S&�omÏ�0�x���bM�Ae�5��%����N���|���T7�6��tT8/�LS�!�ew;&��?Z�P���=�N_i(��~��*�W/� F�\©N�1�*�g@,�9OVZ{X�$v�dQ�x�(�mLΰ�P���8K�wM�f1�B�G3�*��(�3��ڄ⎔���R�PΕz����K�2�p{xV8"u1�G~h�Ҙ���T�jn�s�������2&eք��}��FG��3G��c��̘�epR�a3�������Cg�4�F�n�z���B��$x�)tt�2/;\[�S��E_"V*W�Ȩ������rC��}!�D�sT��+�
�e���b�ه��KQ䓓�u �_bt���X��1< �2EP/��1z�p6��=ze���#�|�?�3���ޫ㬟�g�~Ȇ,��j+*���nw��ʟ��
�O��V���8�G��� ?�u�~�8d�}*��π��q%r�ق����W�\�rS��w��_�����s��]WL�P;�S�M#��e1�g��=Zj���I�7��V��v���N���S[�r׆� ϲ���Ma3�hɱO}�UD����J�"ETD�o�����:@{����QU؄� Y����[���ħ�у���?񹶹�޼����ª�0�絅'f.�|����q2����>B�.�y�\A$�o��~U��I���c�(��c�7�����r��=A���;����A�&6�#.�F6;i�O���c~� ���9���F�nBא4�;�ݶ�ƲujL�����9�W�5p����h�f]�6�yF:^a_z�͒(�HiL����<:�k��X�[��CS�w����L+�j��ra,��j��D%F�5 �s�ODFɪ���L$�͋ �T�{߬����s��TdLrX �S�zf������vO��ʳMV���8>��z���"�{���F3�����;a�,ݔ`T+��)D��+�v��:�՗bUp	:�Z��?��G�h?��ڊ#�z�x���q�l�J`��ƪJE.�� �,n2�H�Q�-hPTW���R����q׊�8��Yhie�L�:�7C�p	/�`�= �1�P�3�Gv����4N?�*�3�f�l�V7����D5�3ȵ�� Z6&�S� �[U�e�Aǡ</��p�Z��:����gΚ�Y��H_3м���]��C�'<�Lz�q����M���	�7iT�$
�G�(=_S\K�yJ�s��=����8u! ��tv�K!���/z�p&�2@��,_o�J�$8���_�'�nR�	��G�}�j&0VēN}3�4z|bǊ��x�_!m盠"���9��A6Z�~_�gV;�[� A|��m��������M�8�9\�����,��P���R}�L '����Kj�����v!rI�C� �����V�jth�r�r�o��݈g�?h$�"Z��B�/G�G�2�ԏ|���;�|�v��3R��rs7l�ϸ:VJ
n3� %eU�"�G���-sAHi��:�4$�4*��bH�N,a>~M:%|�tB��L��a�����>"ap5��D
���r���So�M%���h�W�Eh���w�a�8M�A $D�ν��`j6���K��NE\8Z��V�l��I�����p�n�?9��T+׶L!�jh���T�:�Y4n>���g�T`^+
�Xx��w�������Z�]8����Z�ʱȲ�,Z�@A=��pbrW�����0�j�w�;w&K)=�-7�3�2G�����=u��">Y�vq�Z]|�8L�7�����Y�❱q�����y��ࡈ�����bX$'�����I�V�O*:�OT̟�n�S�&�=����T��Ѽu�V��,���yA LI��:�&X�����w',���ۤu<���J�J�F��*L�#���bgesA�;��B��k�O3�**�gR�zNoWD5���r���C
�Y���r�z�o�)��9�\���n-�����$h\��R�Ս�c՝����B�"�';�cnzܪr�\'%!�m���,%n��7�@p�)�>,��G��YҺR�RL�	~z���R1�8xi��ޅÐ���E�D��~���/ʹs{�KM
�������<�R�c�l���Z9o�(�&
]a6�`YNe����CO��s���]�Lԗ���[���Z�"�4�[�:[}8�C*�Gy+�Ar�k*U_h}q�ɛ�8�2d���Ɓ�xz��=۪i�_'���Ԛ���@$U���R�|6^ma�y�B69�z�l+�2{~��k���q�Bhܥ��T�"�Y��erY��X1��ϒ=��h��c�AD��(/�|�v��N����kp�%HB��}^(&�����E��Tn�3��ǶS����&2�D5�K��\�awd�5Hn8��YZ��������"��]UY�ov�D=s%�e_�ye�:�A��ӱ0M��ِ�C2B���uĚj͔OZq+�����L� f��8+�y�ʣ:�[�ֆ��ϡ��|�_�l>���N�� ��V6[�B7�� �D�>q=��u�Aʝuݎ ����H�l��nȏ�(a�ᅺ9:u0#�h a��K�q�8��w�%�89�p[��
���
���,d{���*��c�.���J�Q����G���T�h���Bm��z�F�����,� ��x ��āH���,WH쬵~|��>l��`llVI'�^�6������Z�	?jM�(yi��r�#@I~�"�Č����L6Pt�1��:	=u7D{x}s�MM�	�Q.�O������t���p�f�W�G�����i$�"2�'���3��mB\�p[�oX�7�9�L&Z��ԉ�|;+�Y���4�.����i�P�Z�W!d��خ�u�,����m49����F3 r�I]�ا�K`g��Ǽ�À�d�6��!Jo�*yo������
�{mR��2�8���?�Iцx����\o<�+��ܩ���#�������u��5�z��%$|�X��H�7���7[���!kY���5��(,��l�'ץ�&P*pzfd�N��I�ڜ:S�����W£�`�=?)���^�49ˡ�c#/��0��x _PD��z���UN�4%�{�-L���6#^i���z�j�2Rz����W�t�wB�?���������!)+>�d9E�>tE�{���+^���'^uJ�G�B]��"�f���yBn��h��kJ����5^��e �"��|)(;�.0W����2tH�k	�K[�Ks����1�ܡ�,�=׭�	�P�Ǚ�q�C����/��f-�\�jZ���o9�Hcu@b. �'<5SD�	�5}Zk�.���o	�^��G����e'>�S1�8�L����sD5�c���q�o�e`�%d丌��{��Gj��Ӄ�j2ǻ�BC�^e����]��6(�O��f籗c�aѭV���`����|���m�����i�uq�vv�9� �Lts����&�QVE|tm�`a��@&���a��tP���'U�R�DO�U�c�81|%<�GT��$�b�;��J>%�+C!2�����be(��)���*h��:ϡWHs�L���Xk�?��΢F9Qi�iՃ�b`h�g���a�6�w��"Ǒ�L����d��ԏQ�.yz�/ɝ` �l�����)�����2�?�psO��s��7掙i�?�O�`���g,t�iC�dҟ*�F���s��H�{�$jp/TJ& Bg8�q�8��|]&�Y�*
Ч����T���\tHx"Iܥw��8�-`m�gtcjM_=��K�tc=A��h�h^�n�8��t9�v����֟T���̈́Z�A-���=>�+�\;[֖�-��!�S��1��sCgS�u�0%��=��� � �0_�@g�Rժd�#-C�'1P2U!����\���Ы���R22�Z��Fj��z��=B;�0�s����A�A>�R��~�f�?�\�����I�p�{ݍC��h���^ 5 �QdmW��ul7��.��I`����I�Q�ExP�ḏ��*�,!�R,"M@�:���z5�u�r�TK�����YOoB�G1��Z��-���b8o׿�j��)8���#���~��@X��E֢!�0M'��p��\�㡯{�'�\�3;�����?s��,�'c�2W��~�{�54��$Lj����i痺�v(+^D����Լ�WU'�r��N��U�pz�`��4�ԎNi���?	�2۔����A$�SK�h�|)<���6�r����n=��cpX[��[Y!�O[W�G�����b�o�|�����  ܪ$L����զ��J�nK"��6�=���?����b�{8q'<�L��:Z��R���'�,�7w��ײ��Ձ�zf�y�e��M)�Z�)�����"���MU�2Q�� . ����f�/mǱF������9�z��P�W����r���]�@��2$M����E!σ�~ � �>3��kb�����Y;3����?n���]�
�=t�跚~��W�\gT�|���"$�6K��c��*�?�F�mQ��.#~S=��r�歍,�+�D��z�6͏�o�Qiѐ�dr���<�e�G��L?0�Ш��k�r���x&��~�f�" �L�~]�XB��K$6��2�������̈́�H�u��݋����Zd���7"�C)0�z7S������P�D�?ȋ�:�Β�g��&I������I���o��2�.i1������.o/�;0�O����E�<������c�,�j;��'���"TA �؀+�,��e{f��ޱ�sl�B��,;�U�5�̳���G�֖�%}0/����()�y��&�G�]�f��X�|��u��[Wp�m�jjd�!�+_ 9�\�cK�0|l7J��z+�F��Ii��=����-�ւa��jQ/@~��_y�k�M;(���/�J�]?6ޝ�� ԧ|w���2X�įt�]��b5��FI,��4=�X�;��!$���[��n%�XN�����sʱ�cY,��F^��y�9�����%���W]���-MS�w���GVT�B�݆q�"c6n�򓙊Y�sS��zN)eBg�r��L�� ��t춤������P5&,��~��9ˇ���%[��`��ã�$!yT�oylJ��n�&�p�S��X�O��B}�a�c�yK�Hb�NOq�#x�k��ゖ[�,�{�r&�e��[���r��F�(V�[���Y=�d������eD̰ϫ�A&@2���N�_�҃��F�����l�k��_S�Au��4�ڦ㧛�7d�5q��Sz�KWr�ܖG
֬||n��b��.2�W��^������XUP�4#�fc,o�g1�&�%�g�!��*�@�[-�Zdes��0i���	�b) _�l��&n�U�BHP/�]0�e��X�H�˜��ޭZ���m���C�mhL�YP��O)sdpgk��!�B�tW9�/*쨵�r�����/�P�b߅�R:��&Q�v��Y�#A��t^�'����n)}�-���	�"zp�f::ҳq�#���X=���˕��5C����J���ې'g�eu���ܰ��'��6bL����{�4pv=���/2�1��)��Q"O�s��Y�/�6U�@#>��&����<�]Pm���R�&�AR��mS
۫/<9��v�b�?A����M�J��xs�Q\�v����(:�&�I7���CS��Q&DS��|̽��$�lu��f��� ��s�l�����g!������s�9@��ػ>QIx�DC��E��̛jg�6��!�Y��uH�a���=�������)+s��&���:�~��-@C�,��~�����mF�L�ށn�{�{���u��r(5��������X�z��fg�����V�9?�̢������-�5H=�������
-��+�b�x]\��JD�pH��u$�Z�U���ɀ�s7�Կ|�Z�(�`�� �W;�#�9[��T����U
/��L�8^��i�=ߟ$�ه�H[��K_�"��@�c������N�P�P;�'�,PxK.��0M�#�(O��R��<H�C���dr�Dv��(P�*�Te�q3@����H^��g*3��E���R��ZT���/��Ѣ��vLٜMÜ�����?�'�v����
����9{odZ�k��p�v��-�x��x""��
�"Lg�ܞ��g�h,:�ag��cdX�p�_�&�W0�yPL���޵��~�bXf���<Ab�Q��	Q��t��c*���L_��ވq��[2�i[�C/�6w8 �,	O�2���>@����pj�:��V�g� ��#{U[� �����¨Ѳ��3kE.{�M�������`+p�Fb�ПcćB��d�!4���i�&�.��<��3\�R�)��6���ri���C��0�]A�M�!��B~o����9�_�\��|X���2*կ���_M�1r��L��.c>K9��3�CK��x!���|Qm��w ~6�(-��u�gN0�s���H���k��25�<4��� ��{��'�r�$	���N��*L{�4��i·3��{��c�e�>� ��ي��w$����u�5FV;Jr����
���W�!g�����~R��WK�G�K\Pn��3�hy���7J�xW7\7:�XZh&�- ����6d���t<�F�H������ʝac4D��K���%��vD����Ed�l"�og_rJ�_4|����um��u�Cn��4��T(�u�e[�|���GX�E7��<-�I����l�=(�%�}�� �'!�gW����ź&��ZK��Y�S�81X{G�)'�Q�\�iD+a8o1i�WqEQB��5��M���y9�9S�l��Y��(�8*�)��9�c�r�
�v`����(�u%�F���� Έ|��R�$`]�XW�]xw^��3iv.`��t�;N4�MX�{�����LZܘt��P��� ��R�fP��(��G�K8���T��wηhl�(L�'u�Ɵ��a�nߠ�8,'8o>�g癵b�C�Cnģ��]���<��D)�@���`]!�SXkX2�[�e�%�o)#� 7ܨ),�J=��UO��Ha����`1Y2i��C���K��)��Yh���f�Z�����q�L�$mѡZ�r�a��:Q���m�g�����m6��<F��ў�Q��1o�B}�ÀG @�Qp#U�ĳzЎ�7W�?u��wu��\@�s����Ұ&�������\���*���{op;���֣o�;,���	-��^�F�Z5S�A6�O�)�-Xq���m4�q��$|%���Ơ�����Wt�f�A�Jo�.�����绲�xY"�nT;��M:Ug�E�,���6u��\<]��+�,�����w^�T�o+/酕vg�>N*�6�
e�`^�����²&o��'�N��ٶ_��kR���P�b��0-�&/�Y���s|�d*Zn5 i��(/�^����6���sr�b�CY�������i�h!�v�A�X�'#��]7O���d�J�e���
K���#U��]cql�dH1E�e��'R�+��=�轘����)����ʮo�^�If�c΢
�<�(�6C ���f�]��vC��;�\Q���3Y=x��4G&A��EJ��_������Ʒ��Ob.|V�����m-"�o�$���%��v2��ʦjj��W|���z��64�$�Vv��WosG߀0���/}�
H3�ƾ��B���ɇ�g���-��+FAPc8ɽ��b�=~�:oA(c���L .M5&�"��s��S���} Z⥌�/BR�Ez�nQ�]X��.�{:JE��̑�(�9�z��@T�$�W�y֋�o�N�w�m�q͵���Kc4��1t��C�D��޾�Lr-K�k̛��P�Ю��6v�Շl�8￢� �6��z�QX�c����3~��5<�����H�4O���^_q](s��۞�mmv��t��_�Z��rEc>�6=�D���N�ƌk]�Ia!m�^\|�Z��>κ�yX��+�N?�l�r���}����M/G��C��/���˸	)�\�$D+w���J4�?\o�N�풇���7��%P���-P#o���"4y~ർ�(�mq�G
q�K[�ZK<�Rh���E��`�#�m�P_>9N_ /e0��c������XY�Ҙ�%���[]5yN �  ���z�v���æY�t�Ɋ���(*#�#��αt��b��1@����� [P
,n�$��8c�t|$��		l�#����Ы�ϙ���H�b�µt�'�D1�1j;��QD@Xf1���Ӓ-�ۃC�M�3��)ُ�d�Aw��2� ��Q����U�L���0������Q��T,��i���t
��I�|U,6��F7��jv���~EF�W��1(�~/�~�ۑ-��Bw4���0����U�4�n+�4���C�S��6��f����g�.z�+-���(������}A����Q)�i!-K51��ǟR~����Z��f�/6T۱9g�E��Sv 5��p��"����~L���"MY�����yФYOyy�Wf��s4f�M|Y1?��*��װ)4O�2��HC�w�mڒ7U��ֶT6A�W�<��y
F�lʈX8ԫ���.LA����H%�!Y~]\`H.?4Tԣm���e ��dD5�d��{�;ҚP&�*�:��֩�X	�`�EP��l�K��64� 
��x{3bυ��>����k�9t9���˱�e�?�/~ۿC����z#�~�	��;e�ׂJ��7�c>�OH��k��f$k������(�J�5��GɅ����30n��E�����{ e5Ƌ8Yѹ"���X4;1�����8^2�UJơ'�H��A��wN!,<�|�k���k�����Ր�`��{��vwDği�հb�!Tҕ�����%�AVQeV�"C�M]d��;$)�Y����/Z��ᓷ�.���П�0ڎCËC9��4J�m��!�q0�����o!���C n�tX��6�>*GM4�3����o����OZ����	�~ĳAsܖQ���{G���yX�x��u��`��\U7<3	ځSk�S�UZ|�77�ˤRnA��l���r�ѳ�������[�5���k������J5���&� ��B6c���c���k���}���m�:G��ǖ��(�U�L����R��Ź��������ظ K���]���gUۉ۸�A�s�|�oQ��q#�i���%��b��<��.A�z��T9�0N�\����GY����B���/�%d���a��Ҁ����~g��ҹ�v��$f>�&y�󃨝����Z�(u�"P��z��
p��G��)�>;��"��u$(Lk�����}K�#�����-.,"�5�_(��Q�𸥋�K^�#u���W)�P��<�Nr��@�&�y0���q�'{�3�KΟ��O"���j�a����I4N$�߮�*#������f��Q5�G��nyv�}0,Vc��p �e��7��W�$���T�+%&j�}����e�Q��OS�
�Y�$��d:��"&+�]�_�[y�����Q	$��ˏ��,Gx'+�"�*��'m�o���Q}s�3�ґ�>8�k���O��d�-O���C>��,1�`��=�Ǝ�m�%�ڜ����4���粺��g^�+���E�`�5Vp�ߢ{yP�{�c+�J�z��bNug�P�y�@O�e����mY�t}_V�k$��R�z,�tx�Ե�дLpq#��y���(vCS�~u;�n�G���f�w&@ ��A3/�"lۉ�ro/��!��"́�ueD�e-xj��T��f�g �����5��N��
�Le�d�Z+���+�k;�.�Βj֯�f�[������9�x���Ӑ��	�[W��S������ԷObP+Hd�/E�֟&X���@7v�bf�'g�fj�����LOœj��w/��%�~0�N�Ț��&��� �5ԇ$�5Cs����:�JS�8A_�B�M�{-�b��kpH��2+�t��Ċ��
_��9p�~�`&Okڧ�/����g����(17�TYTF��Ӂ:C�'"Or����\�\V^�:����X"�mFf}⛴�0, �l��]𰰂����;�߉ �>����}��=%:�D�zg���pԾI�UV��Йy�g���g\\s������!U��~/	�)7��<�ڝ��7#��7q�Pa͔��rm��V���j�v��2"��ܛ�Nܚ�К.gI2��yݻxb%7����uֲ�T[��k��*>m`&�;�OFi>�08��_�!�<��@�L[w��Ɣ7�N�U�°��d<a��Xc�$̿�3���[k�aLG�a��j����%�F�k�wP/n� �b���U\�
**��|���¿?&nf:�!��^:��Ħ-�1����qN�\ȇ�5p�;�,k��R����EfNZ�3~~?Ho+-���Z��y9^�6�
U� �m��.��5�&CeQ�N�(b�;�Y��w��	s�CD�J��Q0e(,���)��j�w�T��Yo��KO���7]2���G��e��b���$�ef�0�j{2@���ㅢ��e"�C����)|�YL���"�͞�)Q6�X�`������Ff`X����$��;����M3.�t�I��~_�s��c#d�Æ+ۥq17&N��X��4��ڟ��w#��Q^~����к!g�3T���X��A:�3	�&�n��a����wD�w9i�"אx<Se�޳���`p��$[d��v��p�.8� �b�oU�-��]m���LƜQ�l�4�"})U����K�n�P�|���������1�e��[g�$?ǂ����@��4O�����6w,�)�k�]0��� ���W۪g�����Ʋ�(��.q��}x�sF�A�1DS���9��j�T�����u8%w++���r£ے<�c�\��_귗�؝⥿�^֙ߘ�$J�q��[��^�ӔZZR��fԵZ�&�t����A�I���3����4K���k�����ixU�}8��c����j�r��-�Vp�Þ5�!�F���duLm/���.�"�Ï:����.�'�>��u�t�����j�JIo�B���_y|�;�`��.Zw��9x}�c��L��W����ٍ����Yv�34��)�E�~���%�ɯ�h+�&Ês������c1��`̅>b��1�W{�vR����g�]-�l�U]%G�_|�R\{+�3�(��N6Li?�;���#Bq�l���
�m<��<`%Ơ��õp���ŀQ�����M�(���n>��P�	��݀�p#��0ͫ�A�Q%G���)D����Z|Pՙ�}7��,�Mq��/<��S�
��w�����W9o�H�[ߐ�uh��J�J�GVk��/�T����4������Y[�w�	8�CJ�*�0z�L���,���
C��ݻ�;�����䭨�tBi��dl���.G�L"Z���ݹ@�v��4��ҁ����̃<!((Dnv&/QV�}|/�u%p��5�
	�3W�t4�o�E@S4�c��W�RC2QL�A��@��!��i�1��6᭛�7N��?�\P�Aj�v�uw�����d*� ��p�Mk�˨Gv���*EV�|)>�ن��� )�1�OgK-�Х�*)WϘo#.��A�>��`��k*��ܟ�k6 (Z�|����l�0�מ1��j�m�e�=U\��g_�W+ӓ��q+>��תD�AU�EgҜQ��k��5t�#%�XO��q�3d+�]$4"�0Z�{�rlq�ϊx��M2,����tb�_b��*�8�r[��MO��J��K(�Ʈ���{�b�Al�?�iM�����n�Xg��)�3&UA0���2�6Ґ����Wbw[�ݐ����~�v\^�9��:Z�b=��,���W����ʍ��#�r�9q���?n[>rl(ps��T�+���.�.����Q�)�c�v�ti�&v�sЋŤ!t�gcL��+j\@�7��Y�b�#�-Fp��Н-l�4��}f�D~�s8�N�� ��R�c�ywד�20�Ԁ�4�Z.�G�C*\_�ԕ 
_|������s���\�;������r��8����g�Mt�G�<G/��s��~M3j\>D�M�I1�b,'�%��|��Vk��֎/�򹞩��#���,��`%BD��]�v���!G�6� �t������6���0��Yz���h�Ν��������ۓ��D̷1���깪�0�`���:�)JÑҾ�
��mU�kǹv��Ji�7�z�����z��榑�Sm�77Fy ;�sJM�*b|
��2���P*C
舥��3�=4�|�Ǭx�c>�����jWE�nߌ�����oٗ�o��J��U�7��XP�2�=��ߓ�fG�}Y�YEj1<V
��+nwI��vB���Ka[~xڳw�<�4�J|�U�F6�C��l��K+�]���3�Q�h�����K�
^���!ᄟ�7��R���ڽ�b��y�D�cS��<�2L�%�F~v2�"#��~���\[����,L�y�\)�E��O��x߁�"�t$e)a����&��yW�m�!Y�(s��ҳgn&��v�D�%�'�B���=��v˼��ewP��p_xe�<�� ʱ�(�����g��')I�ZXIt��B{58��}r�^�m�-�D0{왉)CԹ뭑b���V�^��ڭ���+�[�)�
0���F�Z�����	r��������{6�I�$S��ʻ{�,�F��w����o�fΒ>`fQB��uҎrB� A!���R_g��6�����y�=��6�r�[��M��%Ř����Nxp�ɪ��J7<�����hߗ�*Frl>a�ű�^QoL��wÜ�����\T� F�{�.iI쬥i-��^�Y�p�p1���3pV�K!%��Xx�T����rg�g+���U�Z����1��bpQ7�+\��<�|*���z�F�V�ЀA/%G��b�%c��Pw6���W���~۞&�:�qu����{���?=g�]<D���.+������&ZƄ�qD�U��w禩�����$t�?N��SG�30ID7|�w�MM�쾡���%{z$���X�8�n��
��v�֤����=�db�U�e�x
��D���Nݯ+M�����Vǡ����	r�K-���o�I���n�r��}rV��0V.�:�giW����Kh��V1���X���'�G�܎ԛ�(���N*���I,5���Q�G���y�XiFO@��j��Dވg��t!jz{۳�υ�����qp��(�[(i	��h�1����a�hDS�e���V��Gsu���*(�V�n���1$~T[�
�[����ڳt+9�Y#a�ӧ$�c�[���d����%q��02�����^^�8Xm�R�պ�����yԛ�������1z|t�7�KhE�cz�V;@��������,�-#�\��J~d��;��(�b.ǫ��{kUKy���e�صSױf�2t�h7n�d��8�-BOos���q�R�8�U�u�M8�,��q���~�ܠغs��o�f�)�[�z"`��}��@)����р�k�>� �c�'L,�$_l2 ~ѝ���Ϲ�Df5�����D��pZ���q� �5>!��^��K�h����Hl��]Ñ������vv	��"����P�X�}��YΉ���Y�ׯ��!��	ӆ�5V���6.G�z��!��i����؝ɫ�g�M��^"��ii'�ܯ$S��n���������vb?�}�pVc���A����!��h����kMc���*�5΋�wti��*&<��iVN�7F�ʩ�^���?ٺ�4�d�sI���9{��d�3j��4"�#����9���~ibahP���efv�.IH�'�q�����N��s�ko��6LU�w�� �H�,�q�coR�>��������%
����XP�&�^F��$L��8ղύ ਅE������O�5�,��1F����m,{yk���] �.Z�~��dxF�����1�5;�H�'�dO��q�m�wysr_��%�&�J����9�z�´rw��OsRUZgl�� �ߝhzt|�u���g�z��C�� �mID��U+���|!bOP#7�l���)��~�a�s�b=��<q����t<p��x�9�d��4߯ n�V�]����m�]��6����ӽ�
�4y�L��@�+�]�U���'.�~�-��!-��US
�iV@���R<�pɌ�4(�<�w�iL=�cU"B#,��ݢ2E}_�PC�N�]V҂�[�)ÿ�	�--��~b)����Z�n�|�Չ!xT�{i�h��3��E��3�_�J�����^�F�Tڬ��u�������PG���2�vɉ��f�"��RČ3�X*x	)���jXyXr^���5IX�yס�����8�/�hbQ��Go���i5ۣw����} �1� ��%��Z/~������Y~DXCR��S��z�H��"������a�<,H�V��.����*`at1�nI���~��~�@�(5:8 ���<��I�3����7�py�U
�4Fǚ�H�np��>��-���(cE�#,!
���]��L��i���QL���~=?���k�;»h�Y�4��Ϗ���7�*���&��t���Z�r�`��4f��,$ZD�C�HxKi]yQ��-"q}�ծ�t" �*"���v(�f���
>�l%!le�G&�zcXwX�u����ɜDURO��٤��1�n� $�?aà(�?���T��ܥ6�	-��K"?�b��l�.�_�*�P�O�~�4b_jx��h"[�W=��Oп�s��c
.WQ��|���}F2����!��`������!xf���:��pb��!��띏�1�����8��A����:�:S!�a���s�D����N	%�Q�S�*s"�ķ����[��`�P1��0�>8V�ˍ�?1�s��K�Z�����Sg� �&�y�K-r#��?V�L�Nu����C�.\���=Ӷ�f�]�����<Z"��V�䰧/f@��Qx�V+򭾑W��Ȋ��^�X�Gb���h���8�A@��ҏVE�薾�����C׃��(�S�Ea�'?�x�ry�2�G�;h�A����Ր���������د`�ѵ�x�;�^e���ov^�d���������A�z[f�"+�q�d �|v0Ue�\7��A��R���:�U-���ժ��gm@�F�Ϡ�P�_��CB�8�]L���G��:�0�������r����y�,�^饣�ݯ>����)U��Ҋ0�R�{��&y,��S����_��˾���<����0��_�� �Px�-�����GFZN��j4��QʚOF�k/")}R|	哠���vI<���<*{Z?S�)� ĺ���aG�����6Ӭ�e��e��rx�|?L��I�촸�����-��F���>�Y�b�ƹ�l���5���ր��H�\�����/>x��t�Ϝ<o�����e�A�5���4Ü'�b-G=}�q�x�[����a^Q�R�LԳ���I_>�Ѫ�A�� �*��0�Pt}�����9����21A2d��p�ǋpd'x��+���M!g��S�x	�+���{���@YH���S���8k�,��_,�� �8W�U{���8O���n��u��?�v��x@��OTX� �TοW[���s(�䮸��"w��)%Z��;���$v�{Ň.
�KH��W�dώ��d�ͥX�D�0��Ks��`1̭�."(E�W��\P8r�?�����/ĺċԾ�R�HN�*��pguZ"JPaN��M}%����P��#�4��a�Dp��)z8�-b.a�<�=�s���r[l�8i���(ks#b�p8N�Cr�ˈ��5�'d�5.]���Ζ���s�m3Pbvh�V1��
�a���pP��}h$�2�9`�Y�AZ�]�Ðb�� �#t�vXux/��pX�B esH�IJ����E��6e��LWG�����]Z�����%�ZVX��ɷ���Bo���	W��U�t���TGNT�q���zLX��t���H)-�g�(3���3��j��;�jA�x��r��'L�X�����t��YE�� pr��	�6D[����L�q��dY͸G����?�� \+,v(iw�8.� ,@�ۡ��e��d�`���B0��񔛙_/�{�Z��N"�_�l�J>���9+Aa�i^k�#�"'�u�U�s���/͑�Ɨ�"�*�j� e�~thAO���W���Y?|�#Q��������ʿ��x�Exa^��tq�J�crS�ؚg��n������Z$�`�h�u�-O=��W��e(�pGl?���M��-4��E78��.2y���}MF�h���\���=nD�%�! ��T�'�9`=Kw]���2�����X�ӚG���BJ�T!�"����o8ȋKb�ϧ�Ӿ�[���^,�uY��K̦�Ð��� �"rM}NY[��L���2T�!�������Sl��8���5�c�������1do��;��{>G��9�ެ���J���X�P��X���m�"����x��}��U"��'\��e�k{��z��uL<	XAX"g��x���4GY�֝�K�<˂���kOnY��Ё��'�[[�&@-�r#�9����G'���3�uJ�Yy6�D �~Ǯ�#�I\(�9,�n
q�	.ﶫ$5��l,	ʇ �d�)��q�S6� �ӹ�,k�n��.��h��5�Agzp�R[�U��@(MRG*'r��8D����mSg��%nn-F"���L��hZe��P�o�%b'&V�:��v�D�{5��s��e��{���C�i�nl[sЭ����^�*���&�0@�����nf�� �o �:}+��;���꫆`��"�IİӣB��Ur`�������k,d�5صCk�"&��=��	F��6X�b@���S灶�*W��$O1m]�u�W�`��b\CA"�7� L�QL�)YB.Εj������PP��^�ՙ}!��w���=bL��-R�	A�֣0�B,&�kW*X�Ļ�0 -�9�;����!�@�^�7ܾ�?q\������MtA.n
T1+�v�B��6��;HTF��\��"��l?��?�ip���,���n���(ި��ǃ<����ƙ�ÂW ����~���3�P�:���}i���@
H�1��|lO]!���y~Wp^���%v~��/XO<���8��T?�d~25
5����S2k�'���Q��I>/v��+90�� K��䞾��-�e�P�	�a19�."9��z3�b
$���t�,�#wR�R�kz=a��ղMC��UѼ�����*��?aQ���6qhQN+O�{�`�(�� yyH�{U��a�r���.��@薚�e��y1����=ҍ(K����Y��9��
���E U�݅}�$6��V�H�>祁!9�(���]3^l#��{T��J�4�&4�]�$\a�EKcd�T矊�{9�
$E�5�-���[BH����Mu�ve�|�����Fȉ{��BOx󡼑�\XM�+_,�A]8�@xz6��5�]Kl��]�ZNƞ��"=�Zc���[�_���{�u������E�2�����;aH"�;�a�.�7�6
�]��B5PР����J�B����4�IƳ��fuh5D�ep�E�js�ĲHUq���s�y�
8���h�7�?���%^�L��/�&�㔩�q4s������AF��p^E޽�����D��g�*��F�HNؽ\5��Aɝt�.��/���lL�/Y�}Nf�	Bn�y�>K"t'�1�c4�܃)2~	�#,s�A�և�i��&�VxP����K=!;)�L"�B7?�C	����9�ň�M�-�\�0����wɼ�C��s�AEa�i�X!eq��G���	�ݧۓf�Tbm���Hbt�'G�iYU�ɕ��i����U���p岖|H������RE
���$�fWMRh��T��g/�߸|��z���mB���+Íᒙ���*꿀�J�aA(�^Õ�i.$u��~�ьvi����<omͮ��L���x$��-Z���p�'��v�2uU
��^�g�B\������,�7��W��q���i�AҳVd�����ACI����O��UZ���JE�k���l���*��f�H$��(�l�2��D̫��E�����c0Eј��y|G�ە��6��������D���J��e���$:Fc�(��a�q��q�܌E|vw��T`qp_��ulg�FN���bP~&ы�&���1dXl�.4E[~^ilvP�TH�JЇ��shWZ�`�4^�h��L����{C�Ѯ	��:B#��?<Q��x����p ���Q[n�/�	��Vgs��������WZ��+ρ6Es���X"F�+�V�Z7#FsT��~;�l�}��TC[�$�M1�r6c �������5N��Զ ���3���ö��58R<i%drM��0Ҏ)�2B/��[�je�ɲB��A���"���2al\�����嗃P�8��^���|�������(�
���#������c_
��+Oҧ]MZ%O��\�U,7*4��g�5AT�y��.x�314.��|V " �s��s�D�����YHX�h�;��v��Kh�G���#Q�5�+�<�E��e����+���
�\�����w�����0c�FH^�ctH���V*����{O�kdK�i��^�pA�FCU�}��� �v{���8�'h(�ԍ<@>!1HC �Ά̙��̾�Nt�Ü��*�����h'x���M+X���=Y��x��g�ϛ��ʸFɛm0X�,g�?е���\�j��h�(����AqH������H^Vй,�y>�nŪ�v`��}���2$揑�o%U���Pn�B�y���u�V2W�ޗ�����J���� �(���",f�]n�5"����N�q|��Tl.�3��I&��Qf������"�x6os�o�Դ��4�[�\o(,��>�6w�ǿ��w�J/�)�R�v�7��ei�Aӝ����v�)�\k~�ָĈ'�K�H|���9�ߴ����<����Ve�-J�A<M�V����f��.������I�����-��}t7\c+ͭ��v�(2�����2Н�!K�=s�l��s��_��/��w�lc�����F���|��]�nto�H�Vk%��B�}�� ��V߀&�sU�l��T�;Ie(��Q����J�S��7o�n���<���:������c�>� �N����s�iu@!����ws��fzȯ��?N��O����f��?��J~�K�MMh��T������8��5�aR��lE����Dɤ���NT��u.��"'�h�M�cG�s�K���췮5'ֻH��$t]���U��]X�k��x�2#���Ay0��U��4�Y����Y$s���um�烊}���]��I�#J��ٴ��#�����F�#�.x��a��^h#)1=>�;���=A�x3Ƈ��폸�0p}$���d|�wvZ���^�n��s��6��.0�8z�_h�#�D��'1@�0�-��,|�	�*L��
8+���sR��ݍG�H�80���-���ၽ��s�VҨ�`oydw̝F�qo,}`�:a~)�>���K�N��I�<6 j����n�y�j�ɏ��G[ h:���g��g�uJݯJ^���v�����n�Ga�w.*0(i|^��q^�p�����7��N��wJ8�D̅}�H�ӱe��n�ܣ��J����Y�������B�^"����+ '��Y�ͱ-��莳u�ih��]ڷ>Y]w���!"N&���A�~O�\r�3��F{������0$a)����#e�ޫ�A���� h�'�V,�ּsv	�(���66��"�l5㹔�Z���tyM?�E��P�S�Bq�v�ī"�_F{X���:r��$���!۞��q��0tЪߛ6����V��Axl�(X����9�H�7k�:���[Z�.�hSh�/(Ã��8(+H�m3nFËK�^�~�f}�Kk7�d=̯eb�Q�{ڿy��>����=,{Bc}�6���1��-eX̠?��<��|vX��G@���nz��K��� ���dz��!$���H`r�mǣ`���#S܋�G�b���n���%/l�!���)�{4sx����ω�/Cl�:,N�5^}��@x­�8�ߤ��m<}	9٫�4���ɿ�5ng,�ӎa�F�O���Kf1r�g��:��/=Wbpdۇ�2�y�|��hBr�:|��?NI� q��,Oo���L�1��x�z���<�e�3VY��?F��	/N�P4s�J��L��[AB����ƓȮ���=w�K��$���H���������nJ�g���Ts�[XR\��bϚs���8WW@c�-+Oi�E�#vO����֑t�������5�������!��L��c���8y��I$��dO�i�&���6w��^j�tпjcK�!?/�Qm��CMD�9�/���f�89���3*����Lɮk7����F)��D䋔"�z���ܵkPl�/v�mZP'�^#���sס9�?y��o4�"��p��E�'={����[��p�9G����
��T,
ki|�{�����W��ga{�!X�����$��G"������Y����"~�p����� �ai�y��l���w����F\E|épSҺ���QMҎ��!K2�:Ա0F.�y��蚳�S"�4�1)Z~�"b��ϝ>��Q�J1��Ws  V����(�n�RY��9B!���X��cҬ�t6��(��a���,��6��g�~������\�Y�@���uf�f�w��g��p��J�x�'�9S7�{?��%x�t��T��=�,Xo�7ֆ�@��6r��L�����Za�B���惯��Y�]�)�vs��B;�
.2�H��D��R��a8-��x^��C��8����5���Y�4s�8�H]Zv�������������|ů.�W\3b��Lg��#_��N=;f}Ж-������$�~��n������.�@���H!fkHW���F"���#qՊ��A�3��g�V:�͑�u�=|K�2��t�3����� ����Y%�,�z-_̫��(���� �p���b���'�
6q�.:�L���>e��CH_���I*ĂB���C�\�ȕA�a��b�`Gc7m|եa��1z�`�+��<��n����>������ ����G���H�4�J���g5]��^jZ�كp* �����}D�w��;��\�\\G��2�L�H�Xن2���� Vgw����8�B���7��,�X6��h����Vڢ�P�D0��R��'qŜ�e�/tr'{�\Ȓ�4�?��'2L8X��h~�:��0����]��e�ខ�6�k��!�d���3ak��w�+��*�yܑ-Va��\�(��d��M=1_��T	b���ĝ�*��I*� �"b='�/-�'E�}q���2Ѐ%�2���_��B��Z�_�f�B�[K�K��:���2>r(=o!6�	.n����1�
�t5RU
�Tg��B����H����F�%=/�Fy$�xЂG��4��t���>�ޚ��xҬ�I-xBW�m+���=̿��.j[�No�(j��������(�bj��^�Y����
(æ�S��j��
�l�R�A16w�q�& o�1o��+�֞z�x��Ҏ����,Q;ۄ��@��gD�cIw�Z�6�u$) |V�v��
�*�˛B����k�t�[k[U!��F�,m��������š�mD4tդG"o1
Cu7�"�S|��n�h3��R[���2��>�?�*��T{����<�v�� �(�Y��D�N� ��;C�.���΃T!�Y�3AE)&<�x�.ڟx�@gں�
��Q���(�aW������ �@1��|?sc�Ʃ��ԯ�`�##ݓ�S<��'q�I{o�C�KP��P�I�k��T�$�m=Rn�P���X�$����&[_�X�XW��{&:}�Ќf�=>G'�a��d	r�
q��%�_�;�'������ʿi|
>�
�0~���(uב|#�l�cl�].g7���Lw�8=;*C�U��= ��c���_�dY�V���uT/D�Z;��Y�b��� 6nꖜ�9���ertR��` wK;���JG�����t�T���o:�X;�`z� ��/|r����+��=/���F>��7�A2S��V���5����� �Dg�۝Bn�ȹ� 3���IM̑��I*�ǉ���\!d���2n�!2x�^��|���`�Uzf����f�[9ѣn��;�����c��\�� �7���( �Q�Z�wIU�aG�zJm�������*�W,�#5�e��@b�Q��S��j��*�ދNI���䑗;��f����e��e�gzgl�(T���:KqlA�%�f�M��0F ����Z�Ímh���zpuG߄��%�����b>1�����	����d���t�:�s�j���W6�p�q2��JN0�@/�&+Y��_�hR��l��5u�y����-�Ow��h �a�{��*�C%ӥ��K�"�f]Y�p�肬l�F������g��ʂ\��Q6i��E���ΐn�l�%����ܣ����^��0k~��UCN�@������	֝c�+T}���+�i�K�́���%Ҋ��.�:��F�)>!,�%^�R��AN�3� sz�<�,�\�-Z�}��b��Mc5<�6����d"4�VQ|��<D�3�7�Y�j�*㢣0b\���b��
�Ӝ�y Ig��ʯ�=��	�O�t�O��vf��l��4��0A;[�r���ࣵi|��rЁ�!�w@%�\��2?'��V�����LÈvK�����UI�{')�����6��b<I�����0�� �ՌV�6�)A��Պ��Գ�:�0e�U5�^��f���Os�ݢ�e�K��#�*���O��}�����?�G)��K�mM{�׀���8�l���ho���à�Q�ހ�/���k� W~�g����+�r����L�;���ޒ
��쬷�ߚ���� k*��f\�8낔�'-���7�oB���S�	Z�K�����J�Ď�Sq�`��D�X+D���P�L�UD Y����u�6|���a��s�w{��ń����/�P�"m�*-����&/@�t�U<DkO���>��oXT�H���;a���P;ݿ_}܆����:��w.3�N=ޭ�ל����K�Z@kq,��j�LNg(��cH��=�M�{yәS8 R��ԯ�'u�C��5TSe���}n&۞��(7/����l�h�?���m'{�]��Q���/A	Z�̰��������/�]���jh��٦�,��E=�����ƙ� c�w�[Mt����sJ1�����eM�����_�ta)0F{=^?�/`s�Il��xނ���D4���f:�ͬ+�c�>���[-���cI�͈�L`G	�U�m�rsrn1i\Y���V�9�����E��N7Q�e�gP%���g	��pL�	-�a6�"�=���	�[�-�z�I��n�PA[��#�u����0p0yD���|���r���Շ�:����C��"=(A~3r�X�ڪ���:��W��kR��or����r�Ly6H��GQW��������Vy��R�Ƙ`3�u_<�䟦M�X��|Rs��;b<�F����y.�DHE��Pw�m�1�u�:�rPcq4��y��L��w>�p��W�5�)��2q������lG���P8�ଗy�'EC�7� �����������rYC�T�䢍 ;BzzG��N���W:�N�<b��p���+�Gb����q3q���6���	<G�b�W=�q������G0��:P\��t��^) �[���>�G��ѨeDBa���k�E��4M��5+��*���kk�5���hA��k�
�P�~'ه[���
w��.�B:�CŖ�H�;hKV��t��2�TOga�,�����O��D���1l��b��~��mwUGNtX>��t��%�gf���͞ �9#y~���&�"���X)��o�r��ib�t�섪/���k������դ��z��J;'�h	����R�Yu܉���>�k���D���o�'/��i�~`_>z	����@g�x��-�bE����t;�)H���i���nQ(r3��h6�Yu:��G"����oR׽;��KXZ�+��C�I��b�>��c(����o|̟9H[�k#ցgH6�L����콧aEvT�,�Q͓�.Ł-�������E-]�tAM���/�"q�q�97B�Z��:�~��X�:8+�	Y�������a��U����>���S���á�}T耨2H�0���*�I�ɍ!���&���+z�Uw��#�-5��m���?D����d3c����	g��Ϙ?�cĶ����kN�_e>� ��H�i�#`"+��$�Ы�çŸ!���8o�����E~`�7��������*�S��=0�����>u�8��A��cE�4���Wk�zv!��f�b�L��5�1������</��՟:���R]�&
�kP�� � V�䯖I�/�cS�,�f�;P�� �=�v�
�,���
�4�%��y�X�֍#JfR��Q֗U5��.�&�F�S.`����7�5��QƘ��l�2쥝�������'[/2����\���h��*�}����ձ�6�/������T�����C��qÌ�������n������JX���[U��g>��-r�CwP�X�6�*D+��9�#[2,&K��xp^=6.��^ Qs���ar�uzҗ����ch�z�XZ64Z�Q	�k�óهUj�#k��%���y���|���H���K ��$�@�iQm�܏cTU+A�>�r�>�����#��������ڸl%�@�H/a15�������S���.�0��_��[�o��q���iw��V C=%���0N��%�y����}���R[j�������y;[��Zda�dL��0%_D�������d|���JA,	��$��Hm���.3��8+hX�����ls�Q�`�1�����G~)��2������s�c;�����N��N��O�����z�HyGH���^"�)�#\6�[�����n<�Z�O?@��R\�$�}�1��<�����R7�<�%-�,h��������J�%�� [c{X����ث�2|=O���~ۦ6AK��T��.=	�=�h��T�m��u�}�C4�鈉�ܣ�ƕ�'T��Ń�.��Uv��$������c�`8�;����WMwL|����u�7����o�F|KFX��{�C�A��i�aJA��p7�j��4�Й��FH��\ ��.�$w�x>{t��?	�A{�8����JP�i��B�@#7oq��p=�C�&<�!t�Ի�UU�L,���P oz6���1T��u�)/��Ack;w�0��Ձ��c��/�����ѕ[��>)���S��7vȍw�2��TvqߎI�&R��ԅ�4C&��T!�5�2{
��ϫV��ͅ|c��t�?8���"-�$�Z��X-ֺ^��P��\f%�'��t�Z7�6r�n;H|$���ڀ�Yh�sW������Q�����f����K�%7�9�?1@NpG�-�G����=�j�)M�MМL-�H��K��磛��y�=�9�]�I�y�ﲩ1�2�yn�����W?�j���<N��<ڦ���Ԝ�@�r���� !�X_SCg��r�;cP���I���dOYїO�J|$�x`k�Lho�s�x/bA�L�~�l�[��1�����Ҡg��3��>�	�UX���Q�!Di��8+�]�mB�'�,274G��c*��S6����=��; %�٢�L���M�($�`��'[��י=:y|eϊ6��K];
��~����>����$��RA[�u�<Za��I�V���5�7"I�c�#c^J�xǨ{0���t1P��
o��C��c)x�&R�9�bu���rK?8���"m.&��sggb= ��߄��d��;���6_��,�'���"4{��f^�����a��m��R F�?�m�yod�N܀���i��㹱/�Z��@@=]XV ��\�����;'������3�3:e�J�p�YƬΈ����pl�*Q�L��<ʜ�Y�J@*)��ʦB�E��0Ȩ��x��[�R_���E�Z7u�A�z�}]��z+��c���N���DI��Nݱv39W��Կ���/��l;.֧��9��=�^��V�+�T&DЌ���)C6SI�8����+��{���(I��)U{n ��k^^�n��w���SA�vF恩K�HQ�
�%�tkAW̆;o��:U��Z�2���J>pDX_���X^JJ�(��yT�y�-��V]-�hE��;T���x�LRv���|bߵyQ�2	���*�]d��1>���e��n@򁝭�燢�x�ộ��1�+����o� ��46�و$���7Ϸ���~;<�]�k-�Dy��|S�����K�2ƜJ���re_�G����+��㣽I���Q���TBS=�-��
�^]暎X�MK���&ț�#ڋu[
��{�}�%����:t��c��BJ�:�h\�}eGE:}dD�J!�C��S���]a�p/%��R��w��4��y�sP�-6���b���~���'��}��Pp��8����>��",
}���0$�݁>�Z`�tqYe����<`|�2��f��M#�j�ЭI��{��r��C^�d'��}���6�~.͗�A��6�8*���?^����깬c�W)��Q��߇�%�����S�Z)�Qa�Ch*� ��׮X�O��^@������%�{#_��G��Zgo��~��������%jlS]D.��N����"�7��MXm�|>~ƻ˚����o�+�N��`e�΄DkOu�ж?z�+e'|�����Պ�q�LB���ף�0�>�SD�:��T�*���p��}W��U�E�u�	�'ә[�=��(�7���x�ǻ̀�Qp3n`넅A��H�%�1��?�dw���y��z����^���B�Ŀѿ�� D+J��"C;�����\���S�X�aGV ���yT����QF*bB��Z���>�p/�q���x-{?��ω�� �j��} VQ�ٿ�������rР�G�<��6O-�d�)�*�L��m��̯d���5��v��q���_�#K���a*�y(�G����c�e�u��;�Ω�\�F�d�4�!��-�U���Nx�8n���!F�#Rj�Q���@�bX�P]��8Q��=���5Gw���$�}a���؀5?/}�t�!�42�yH)o���ԡ~����(gq'������*��][Ƴ���q�hr�KS^�~Q:��I��Hn�����B|��?��?����X^,%�L����f�i�@4Z�]#��+��mY$	o�Y��Ԟ�м��ƥ���hE��w�3鹖�W����?#���cQ=d���n��D�{��7�X��?�K���R�"V'��]+�V�lm�����A�&Ǜ�����wl�sa����Tib�H¯�hƮҰdQ}%d⢗���SxY�?��i������.7 x�/Y%���=T+��l� �q=f��{,/���Wk7�D�j~'�Iad[�P�eQ�ɞ-얇�o�T���{�h�wc톸q�y���ҭ���4�Q���ԭ\�z`��{Ky��B�Y�� s*��w�pӱL��-��F'�2xb��`Z�_�;��W��A:��ۛ���F�E�4��32������ab{@�˝7�za�J,���`-#��ӝ���WAҶ�M��S�m^^��Cj߫�}.]�S�LbP�6!h�ODV�J�@:���V��N"�� 楴�\B���D�����bU�)/�LM��c�n���Z��+̔.�d`�4�J��k�Q��ǖM���9�\>(PB�X�睍�Ĥ���d�0��_��%/�,�"s���%Ha��>���P��T�Z`�Y���p�/C L����+671�hG�ZY����W2® S����]����q���TV��޶F?c�jX��e�vuҰ.A�]Qz�YI�#�A�-�����g�k�]:���1�g5�/���&��ѡL�n�*��
��DʘZ�l���8�.��F-�w ��Ԙ��qxFA:@�=T�Fj��
.Z9-���ʥ08�ǟ-��6Q��l�B��j����ݳ�������� ŘSݣџ�b��1z���_��q��XHZ���x"�r�GYƦ����.}u	�f=�����c�7�>���)�2�Аp�xm�Jؠ���t)��;[�qB��)C'��H?%{3�Ҭ5����sM6f<d�62�/^�`���C�ȗ�C%�ZH�P�3.�W�1#��)&u-��-S��}��$�L�@�����~����a�c>f�~�钽F2�����C�X��n��kl�ۿY 1G���d�b��"V�j������tdG���w�Q�G0����k>B}��	��F���J�E���*�nρ�4ǹrӆ����\��e��ꎜr���e�jȼ�C�6���M�n���V�f���"��G�qh	�u�P�kxG��H�ӡe��M��d<+�Da�J]�%��5*#ӝ���C_/�%��CG�@�B��R=A����5��J��m�r3��z{.��]�k:����x�g��۪�B.�r˻4�"/c��-W
��U��D[�*b�L����2�'�7��Ad|�%�����*�m�ê�	��	\��b��Mp�7�4�.-��SG	Ԛ*n�UNi�qqwk���PW炧����#�*Q}N���_�����7=0�PIDb���C���d���io�� ��礰�VB$����0�K�ԽC�v�:jn8^:.���y/��<�����_0S�l�6��5bk�a��ыb�|��\����]"���
� �uK]"�%{zz�Avp戓�AķQm1�r���[	y���\Y���k��9�T��e��l5�c�aV	p�Uv����7W�OK�>z�1!P.4.�#�wN@G-S��V:Ђ�v�[#Hˬ��z�&z]Lk؂�!�p��zcٓf��FE/�0�bq[���9��ӄd����x�.��i�����6�P~�3nɖ��s�!��ao�����!��O�������5�$jA����=(�dvH�\j^�,6Aؕ 2n��WX�_gx�l�t�,'�6�W=c ���T���&.��!2�;���X�&��Wy�S����n�/�o�J=�
���P���ps_���� ��,[�tX'�^7���Q��c�[�i�R�A4}2� 1�4n,
K-�b.DB�q)���Kbx6�!��^�y�C��DW��G.PL���`�"���.�t�-k*��/�N#i�G���:��3�(�-E(T��������\*��X֪ټ�I"߮�M��]f�>�DPi�$�i��#�F'WY����X���]m#�o�6���h,zz�9��IS۫腪���+
�4��}�˄>�<�u߽�!+@��	}���Jgi���#��b;`P�@N�@4����T�!	A|����i	
�K�=B��G�fb/�3��rp%�I�>��1hj�/Q�b5&�L�H��8c$�x�%��4�ed����P�/���-���~o0��@��ua�KR=a��[k��PƧiH:�'�O�b�K�KjoN�"V�o�J�Pz�\�w���N"���B+{@孙�����������=O&Rv�'d$�b�4��ҍ(T�]2ߕ��k#�^���b� \�g�<�M�bp����\>�۔j�?��UtJ:9s����*&s\��:�9V���~P��=�'����c�r�������Z�%Dnf_��;�D ���|2�&�����g��-��L�v;q�r��׼�t�;�0,���+�w,t)��O/�,^��Fj��F�?�ۋ�&����z�2I��։��PC:d�s6Bq���L��EE7�ݙ\d�9!Gp���ӛ�`Z�-��W���rԔ���|_��������]��6����\>A�N��!S,�
��E.���Cs*D��.9��kǾGa� O�)�>��rԊj�Dl���fDٓp��M���)�T���f|N!"��?A�jk/n�A�(�x��vV�EF@��J�/��s�QwҰR�ū�q��8h�1/�
���ˉ%~Q�O�e���f���Pi���+^�~��X����n�5P����K��V���yVc�k�!l��u{�{�lk(��=lwd�=$H�Mڬ,v�+�x�ym�����!S�$4m(�T����Y� �nt��LP��F�m͢��r7]yg��wO��FR���ّ^l#�G����So���?q���-��!'=(z:��g�@C�a:�&�麴�r[�������� �X��`��ژg?�#��HG���+��͟�o�ڎ��F���&��^e���v�Ç����2&+�XX�կ�^�C��-�c�N����y܁���R�z�c)��?�("�K�>hT��BSfy���)p�.D�A�yn�*���:שղ�Nh�kr��}�M�qQ���V���Rb[����)�c�Z�(V��a������[��ʦu��	 d��z����m��M8�)S;>8�*6��Ú������R�O@���xvP
��ğ��T�U�L���5�c_�M�^^'�B��w��sJ��K��M�\��I8�Vݜ\A�N8�U4j��)n
̺2,���W� n����_ŝ쏉Ð�w��m�M��x��DY��7pn���]���XZ�I�( ��H�H<��q2�`o����������s9��*L�6�fL</�Ќ��s�$�o�rvq���'���8��љl��=��Mξ�$��5�Q��Yy\+�>�UBVvK'�bQ�`r��;@='<O_�f|ϲ��:�IAu��ؐ8x��%��᫶8��]���P.ytI��	�����y܇s��& ?K�	b�ܹϦr/ ~�\���+�;���?��l)�X9�T��z�)�0luof��ꖭ�6�2].]��	F�V͝a߫����zq��>�����@�VB@C��Y*N�.���q����� �x(ۥ�[��M����}~D�U����z�P�G�M�'�	}K̏��T���SE���T�R�3^0��=��k�8A����`�=۲�?�-���%Æ%t5i0���j�S��0f@�Y`9�fS�2�����j�Ȭ^[x ��%����s?3m�d_*���I� ���z��_Oht�eD���*���+g�.�l��� �;�\E������D��q�4��j����֎ԟ����KV9��Y��|�I-^���A��Ϣ�����U���Tln�*R�FR�6��&6Pe�����é��֜R�Y:�a��͓������&�=V^F�T6���{��hU���_J�rh�[�FR�#�W$����6�"�l6�sR-��L5Qÿ���,9m5(7I�eAw�D\���\�+��/�<�.RS����w�r�������i�UȆ�vؖ�?��	@d�Oj�4�)3׉��� .T��u5��eU���Z����̾�?��`���Z��¢��ðl��{�l"��9��L����@�aY�� �|�?PD�.�\e����� M6E��?�&=�z��{�m���2��������k5"��m�r?���d�!	v҇��#�m8:(0����[*�����Tz�r��o ��'�aj���x�S$��oGh��ķSD�
�?�S��&B�nr$y�-Y���f꒣~]/�W�+9y���1ǑIk�fO�,F����F�d��� A�
�H��f�Sm�d�Dw�hr�0$AR�W��`�����g`r�b������V,U�r�Wܥ�9w �`C���N{�����d�鏻��O�84*Q�.�O�5����Èx�H��˖SbyU�f�q�_}��#�2t+�T�����Q����d�w�}h�ߜ�8ˌ��X�l0B ��r�쒂��%�O�t�]��s�$(J��7����*BO�����NAFb,�y��X�X�#_��L�r�����"�JHv��?�0��b����f.s�6'U����dX&o�'E ���cyb�s!�ګ�f��(�7Bem֡��	5�"��)b��М	�u[Ȭ#�}�6�t��L�X��&��;���f`���Z;�2��ߔ�;����2r�6�z�wƀL#7_I.v�1�s�Ҭ�h�G�8�HY1�fA��O�ͫ�����f�}���e�]�jX9��%k����.��HR��9#=�'y��O��^Vټ���d����\�圃�u�<:(��k��p����Tq�G��~ٿ����L�o�1�H�{�7��0h4��G���!P�D�Ċt��>EgZ�'}�6��EMX�f%��k�ӗ�	ՠS�G1g�l��T�х�%]�Bdş��P� ��;#��96m�Ե��J������l\��	Ӄ�j�$��4�<���Q��^�XC��c{Yg�3!~Ó		L<j�*q�`�"�Rꮆ�k��d�x#�ώ5�	qr��h;悊:����t�*��
�m.v�:���q�ΠW�P�p���Yҡ�t�+$� L�i>���>`��a��|��-2p�vid$��s���խ_��֟1�r+�����ѷ��H����~�20~_�k�ª�1�!�E|k4�&�,DUN�#�]�pٵ��8��4�p����-ב���As𛿺c���������8NHr��/�%���"d��d��Ƿ�Ď�q�b��s^�d�Bٮ��A���nO�Yj�/^���Ep����&��ډ��p�;�ņN2�xW�d��J{s���6m
���zhJ�Sj��m���Xf̑�ރ�B�	0��a�Ӫf9�C�6�P�8I
_�1F<t=�b�0F��� �� M�!�$ҫ���{�9�~-�Yd�|�v�<��(T˯�
�9�Ge{;md�y�p������txNqu����{t6�g% .�5$�Vo�V�*bYH��h+�`�!,㭍:�pş�d�{Fw��2�3�S�n|�d�˵3;���Df���Y]{ �0�E�R� #�/��"0����'"s;�]J���c�׎>��a��Xj�S�u>	#���b�ě���UF 6��0��hզ���?�%�������C�T<С��x6j7\�B���jτ�ǀ�h����ę��3��n%���kl1x�`����<�s�DL���x�=���aA	��B;����F���d��Mz�R���8{�h.МD�m�Cbʫ���~lx��#�K�"����G�wN����������s�A:�I;)�����{����� tt�U�J�c�!�(���2�d�s@SƗ2�Ġ$2̖�I�7Z�e?�;F�$�9h�)u^���A���7�T��0���wDY����W�{�I�S�&"���U[V.�@1��n9���%EP�p=q�nh�w[ _b;4��"=��籮������A5����;�$:ė�m�������0���#T� ���T�������˪{ )y�^��UE��x,���itMB���q�F���F��K���W���L���.�I0oO^��q��S'fD�$����\(}@j�p��5K �S�y��R�e˶_ʩ��K3���y��_*�1�x%�)N��'�#��͕춹�z�en�8-�����{u��l���Y�l?�eY�!cѣ�v�^�>���^���jJ1e�:V����<�J;m"}�5.��8��9!%hq�Ss �y�ο��s��Y��F��փ���#�*��<.Pg��&���Y��
/�1'8��g�'So��ޮ��7��r�������2e���E�����7kۻDֱ��ڝ��Ѡ42Cop��9���0J\��J��;���爖�e����Z���P��H�����m�0�f 2�lt��׷���L�|瓒��h��O)
w�_h26wܖ���hX�4E��Y��D�����8�v1�CEm��U	���D4ӯ�,נ\L�:>P6�N��.]�������a�(���7�Zb,�	n܈��E('#�uD�I��Y1�1�I�BOl�Um*ඈ mp歗�`~6�*j�@'���RѸ���"H��q�k�����[�?�^`}��{�;��Wxb3�߶9��4��\��1v�,�<�u&�Q��SFbn)S�Ȥ��>��ʉ�H��f�~� +&o��갗��k�-c2r��P�u3`;�։I�)�xY�K�w�4���~�!]�R���:��E<FPBUM��W��>�%�4�n�;ۮ�(�s*(C n�@��^���= ��կ"���d�p�\Ij�G�$�S>�-j�&܏8�(�q���s�p?{ .���^ �{{��+�����>Bi�~�Q9�:�5�!�
$��oK���e�S7W�ԋ�jD;4�����-���R<;���ntիb�H���%�QB��W'���J>y,�c���RO9���5h0-Zz����#r'��  ��se�
Z�;늰�)0f�eS�+���0�h�ڰVT��������b���2��œ�"�#�s�Llߚ;#�k�'�����ɩ�2�Ш0����M�:��KnUOUDdu��@g�|�o�Y"�	5���<�h�a/o�^w�U 5�=�o�'G�,~j<5�JM�D��=��p�<nh,7��N��B���o�`�̴��F���%�,����8gAX�_s d俌n[m�(y�?��4j�t����N�o,'��u�f��yL2&>s F���uZ/��g�`nw��}i���Խ�[|����c����vxH.�A�u���'(�N���s�9�Z���?�SV�C��cR���i7������&�/��8l�ш�q9d��a�����A�v�;/�7_E ��&�*8p^��Mn�c�y=V%5��Y���q���sv?��:d���9#T��l^��3V�M�X,��7_!����4g.�<W��fFc��NQ���v����?��O�q�����xX�8�)ؘ��=��|���WMS�-��j���G	� �+��{RG���m���H������:��qRL2��Vۺ�A<�B����e���t�w9��>��PX�]�NB�O���$�!<n�١��/���Ef���~�))͍eW�6u .��Fj�>=D��IOҳb"6�}��뇁�йNf���+cN
Miă���t�3� �`�z��Sm�ca���Z2S���N�,ܾ���x�s�F�w�%-��#ر��cq ��L�<��'d3Q˪Q��Ylf����ϲ����m '�nhn����,�~e�����)�D�Ip���>�[���H�4����c�ϥ&��1��+w�/$��̹����6��aԋ]�"Ţ>T���a�5�VJ����4N�4L��'N~7������n�ҿ��0M}n���-p�!�ǎ���F���Cw��fdE�b~i7H�l{�L�hvedeV����}	��Mt��A0FǦfer����1?�p\óG�:�@i޲&L4�6w�]�)}?_`\L\d���꫍:ELp䧃�d:��chӸW�J
���K�"60��oΩ��cM��폝�t�
8�ِ;[^�CsŘ�{6*�	�4�3���P	�r ���+�J-��&6�,��]�J`�[���ЍjLA��8-!s��������͙�b��1�0X��(ğ��y���f�g�u��w��?Z��GN9B�1�t	I����~�JN��q)1s����'��^�x� ghH5 �Q�@����zV*�(�ē�ʟ�Wľ<�VG�����R�L�,���kE�3�.���'�(x�^u�W�1E������ ���V���)T���$/��eğ�+�b���x�Q����O�8vc�^�:�&1;����[wD��,5��]!��^��X��/`��)�ӌvv����C�Dp�=�[t�?ц��܀�^.�(�G5N����1�9+�����LѲ|���:�K�_	/jUtw�_\�TF��mJ������7to����Ws����M�}죍��ո�����ʢ���a0���O�c����=%�xl�[ ��ߖ�����n�:��t��@�nB��R��3��x�o9��zsY|�h��Z���	Q���uY+s$�5��㧑M�M󄘚n��S�)�iUDoA^�*�n�!�
���/�
R���;n�&:&�� ����.�Q`����8��"��5��h���r�:���O�����̶�$۸�B��L �ǖ�wm���c��8�?q����B'�NY|�������o�_M��%טp���\)e/�=�D�7�w� �+w���O���ĝ��c��e�hM�26ő�܋N�j�R[Ƭ���׮X�WPj�}1��8��YK<��ڙ9���gCNC"�bB���5��g��5f�ŏ��6�)~��\$����r2Nk�T�C�Ab����	E���'�gn���A\n]���,�{����&�Wy���M�<��tK��eǟ ���'^_D^�������
d�J��f���ݭ�܍j�*q]ѐ���(^�qy��V_�ܺ�_�eB�/�2��E���S7�H��}:�LTl�3u2/��A�8@սhxL�-;˷.rX�6ڥ����=�9+il�	�߈R�5�˹d��nH��/�?'� �J�|����oN���R��ݝ S�Nn�Ag�J�@�����kG�d�}�I��v͞����Eq%,�Z��YJ�'�Z!͍��Cv�
ϝ��v�F�B�0�{̡�O,V�>`������|���3EW��f�CM|�א�pƶx���@2� �TD��+�c�ޟ̄���tv6����D�����A��=@�'�.�QeV:%(�f<lMڜ����?p'ze�O�����0�(����m�x�j����J{K��\ЂL��֖G�I����X���j��	6&��ʙ�Ĭ`Ӝ��}�l^pY&g����E���=��ZL��1����R
ua���x=^���N+�zh���Z�s��/��=T((��L�~�n��ٴFh��*�V1��]Q�$�PPxxa�vm%D��򾎸
��i�%+�%VL����$f��h�3�l���0�T���V�$�*x*g�'�l��j�3K��efX x�5JJ Q�>�������!^jbOz���Lv�%�9�T5۪*5پ���(���.p	��\�̹#YN	p�.`��q�]s�^��|�Q�0�"@+�*�M�9ܲڨ����(a�Cm0SӅ�u|���Uو��= �aؑy�y1���U�L��@O�F)HY��B�Xn�_斝�l�[����Z!q�x�:�ډg��&�VfG������I,��J2fC�;����c��J5�� /���K�F�zW�h��0���a��vd*��g2 ���]��*
Y���b�8������:I@��R�;��,9�;o���O�4>�-U@g/;"��X�o(�Ыڑǻ�+�K� gx�����w�&�����|(}3����"�Ғp�N�&�����@�+��p�i�;υӏ��/�C�鄶j -p��'C@.�gZUB�?�1��0QX�ɖ�����lѻ �W3"��?s������daW�*?Bdx.��a~�w���܁�!��͇�Q����f�V��
~7#�+h{Vl�Q�{��q���!'��,u�MPV�H����ŵ��<G�Jp���	?n7� ����%5cM�k5�zzJ����$eCp���w�S�N*��"W%Q���D�Vս�������s�u%g��ם����gZ���Z9a��"����o.U0wC�f���$/#�0��q>�8q��x�3&BM�vqb�;��P-��Cv�4dNsθ���iDK?�S�4!@\-�W��M��M{�>+^~!q{�S��3����Ju���(pA�t��q��@��M���H�"i!A�t麧rxq���)���_�˝�אL�����{�'�VON�/�Ω� c��*G��_6>y��)3�}�.�s�c�ä��rd�#�ȏ����~1����~l�E�o��E����U� �7�8�LW	`
V�_�OA���59i�"��JCԬ黁��&���|`�* �̰��u�xBpms20qQ�����>,waGwG�9�x3T�L��8�R��)����h����H	"��Cū�I�v��8�p-�!E���CO�S`w�(T�W�vBDm��ޣ-7��>��l�j^>��pd��$�7�=��sWZ1'c㉝#���#|֠�ٽ]pj%�k�Y��Y�ab��J|��p��9n��cK�SM[ؘ��qp����	�|1�����_mr�?�}�*A���Y3=�$��$�p7�ɯ���	���-���0,�S�o��Z���L�}T��[ss!��j��P�T\�	B������t��ԽAѪp$�� ��k5�C�A������a>���n&���Hy�5�?�����%@�y��Hz�"D�N2%�R,bD@)���7��+gV��tD�'IWzP1��*����CH�h��kn�>�ԭB9��YE�q���2�i(��QL���`���ZƈT��U��Kؓ���gk�p�����K�R��[`�a�G���A�����2/E'o�8�ڪ{�ϡ`�#��	'*���QS�zo��O������LA�'|�#����6��v% !u�H�Of�^� �ځ-��-�Pp"����7n�Tͨ�+5�k�r*l������v��o��L�Ӌ�����9��$�\|.��a�r:�{�qh嬵��	lJE䤱5��$2�V������֯#�M�����?wq#	s94R�?��k�F�G�����~�� ��Ӳ�W�8�3p��qge�����?�~V�ӹ�����4���A5<X���_�{y:i��똿�Hy��S#�e>�-��8��p�����:�x��z%v��z�5�$}�wK5�<p3Lt��"�'0���jR����?�.�$Z�`a\h_!��Aq�kTy�>!��m�Ɔ b����?<�z�Qo�G�l��� "���9K_}�Kj9Qk�D@���َ��|d��^m
�j`�Z
^�Q����b�a�8��m?���k�����RW�JW���4RFw\eU���(�����r|��l�٥��}NC�^5u���sX�ЂY�7oI{��m=2,�:�y[Ɨ>����OV�+����
�ǳ����Be�������ׂ�:DJ�pp0d_�i��;.��M6?�$Ϟ�*"��,�h։	���An�j���0O�'��	R���U�t��!e6��M�E܁;$�/'t���ٯ,.*�V���j�%M.W)��J���U ���*�r�E�Pe+Ǥ[�ʂ�����bV6C�M@D�^�!)E|a��N�HOr�[l�1��N����[�`��vp�$F|��QEÕ�F�oT�z@3��	�Ih�sz��M^{����cϹC���A�J�a	YQ61���N?�i��`c�?�������c�񜩪9�s��N���d1��t6ѡ08�h�z�6hE���в )���Ч4k�i�+�Y�
q4^�>���}��a,{�Dy��+�ʭ�����g��f��ֱ=�������c�Dk�RQq�S�l�g����c�J)��=�B5S�o�r�pH�>�*iK.�G�2��;a�0t�(��&���_��V�=��>������Hą~a=�Z1��Ķ�mWYF2ä��(GJ�����ZM�.�re�]HO}n�=�(m�=Q�x�Rg�</.<�TY��
��,pEd�{�=��-�9^w�Ji��)J�P��7�+��'}Y>֚t��*�����eW<�#>��r�	��g�I��0]�k�}ѰB0ܭ_oؖ��S�=����v���RS���#k�p��<`����%��+ aK�4}���b��x�q�s�s�+
j��>�`U���3��ڌ�f�g�M���s޹Fp���Q���w�r�@16d�@�3;p��������R��gb��ǣSa�#`��@Ø"�ao��ln��bWFt�uu��?��4�:J%���G�zZ�����N�]R�"�� �gMũ['�&��~��J����S�R����m�*"�L������oL�߅�ⴈQ�@[�͠`��
�HM��r�pA�H���W�f�RO��F>l�i`���ҩ��'iW���L#�$7�7%�C8GM
%�/�gt�L,ʠ��zlGj#�L�L�,gєJ����?/�<6�o��%��,��k���a�E�3R]�#|6IK��P��܊R�^Ђ�:.�Ἇ>S�Y567\��58�����n�F&T��::�맫�TH��� �Xa��C	��e�%}5xXaz�W6��֞nA�]q��i���_�}p<�����71�DG'�7o�X�w���PH�B�{��Jft�Z?B3E�h�\�Ņ�wg��	6���s�`(�6�#��4,�o�jl��(��@K�'˰�D�����j�DR<��T�%-��
����v����)�����ʨ'LÄc+N���z�#}�s L�H�1M՟�m,���7D�M�h����pQ<5rI���a����<�|#���X���˽P*���W[�9)�9 v��qS��N��^hAyV�3K�>�����N����c%����4�^bC����X1�	��/��>�-6ҟ*)�pZ��e�E\+ܝ{�v�s��B�|�ٻ2��;����9o>6_w�*��y9�+$�'���D�Ö������,V�^vTE�G�(=w�G�8c�	�c.�6����/Yu�Z��u:�j����.!:̽�n�H���˿�}�eT��B�$dU�۞W6�D�})'OG���l�*�%yc�%�C��؂[�R�K��(͙����=μ��.UG��g6�a^X,�-��^����(-�{�,�����ҽ2�yI�6��4�<���ا�.<v��BWb˧a�=��w5�_�@$���ʲ�v�-Ը�-�8��#si���" �Z�G��^�{�]�W�{�r~��׉+��bZ�! ��`�Ѩ�4=��nW����I\�sؙ��c�ߍOW*�H�����Pl'?����xHX�|a���tԵNpN6�*�w��ѵ��u�Iv��g������0Ue�K=�r��{kތ�C20&}�`�Ӌ(�N��>����B��3t߄�_�N��B�u���ܲ�x�����J���-^��~�j8,�_qn z,�b`	��X�����v��b.�\ ����@�=QQ�H^̳��
:�n�˷I�S.��l5Y�T�e��i�Yma��r�X���n�
�4��S0c��:��!��t�/
&	�ࣨ�v,-�RR����m�ǹ�o�e-h��Q����Ȫޘ�p+qd�(������Z=�:e�1�j��1pO����F�W3t��
�l�(?C�ww$hs͢����_�ƹ�lᑶ�hC��L���\��Z�`��М-��a���Ňmg��3�6���+�s ;y>��:���N%��W!�6���G���n��F�6S�g��#e5��`jɂ�^�"	�+�0��b_�A�k1�٧����j�٥x�~d�P�M�r�h��lP�g֛��F�x�^�1%�����`>�e�2�Ȇȡ�l�֟	�v1O��4��x �R�*�-�5�Ѯ��?c'��K4�	� Q��t8 5�(�NDuV�4fT_x6��°�������Ǘ�fq��iY�OFe�s�҇���T�!Ҵ�u���|W���8��*�~+*.k*�W���z�z���>�eq��0&
}e)T ��=C�C��>l�z��s�`�Sv|�!6)<�r��蜏(���^x��J�|�:���|�_���Ÿ�g�V���[w��7�*�5�"/WG����%� M��bt����|2HF��Y .U�v��&Z'ߣt�+�X�T��/�[��t�k�q�pxj��i省���Ya�y%l���.*-c(��T}�M����N??&F��$�f��}w&bR�un��l� -yZ��a�0-�%J�N��M���3��D�$r��+��41^F���֙���h�������,����f�(�5Mĕ�%̀�r����=|N�a47L��M �@U�r�z��8|}`��P�}��_v���[_ �?��|,>�YO�?� Ǖ
���<�K=O��-����H,��'2"_bL �@@�������=�<�|r0�r&A��l�F/���3��B�^$	
�,�J������;tO�H��͐�o���s�Ǟ�����o ��F�y�h�)�oCe�C��nbD�!K���%�k�I4�yWzYIaNz����u���!�~�<he��]���aWA�>k��,�YB�I���*|�t0�9�n��9N���5��죡|��7u#�7��4g�kY0����F��+y,�:h�����tkD��{�+��Q28�o@bҫ��#r`�Ky��H���Ů��śB���\�{�3	��k�8~��xy!�x����*ܥC!����ٹGB�?�?�e�t����N��'���D��}��߼�<���
����Ri^0�u����h%7��ФƸ�)���l��������(�b��Kw�ϕf��z��g���6ȷ�\��j��Y����m_�P�M�0�1�-Z%gb0+��3��J��)�,	*��:Vkl�gxe]9��y�L(J2\$��o��N��Y&���S���Da�qj~ w��/Fi7av�3ܳ�w ���O&������U��YYeep"[�ov�����a��8����+y��_���]pE`�>�6��zKuy'�R��C;��S-�i��j����k�g-�K�I����v �J
t0�c�&5�ƁG7T����6�A�V�M5���e���KA�ם"�!2�0����^��{R+�́�����a�3���j��fvv=�ő����{D,���z3V�Njb'��RA�XE�2������*�-D�ip��g�x.��-{n���[\�*�VIp��;;�� p�`4�[��୞������ݏ�}1حVg��u���ҭ���k�zɷ
���8��;hx:�Tw]ɥm����5��z6Ũ�����l�`]@k�n��5�G�1Gy�,��`�-��/$��٠^C�k�CD^�o���c4�#���ܣQ��OOQA�%8�(hPcƾ�m83:��g������y�XvS�q��dδ�*[����d�  `5��R��J�i>W����ऋ��j��`4y>�x�7[���Gُ�L��?�/y�BIΧ�N
e\��/I�r�l���w��6^�a��A�pW{�PP�t5��sG8Hr�C�#<hp��{qG���_��6H�'w���\8Wwnc�����I�n�6�Ҙ��!&��J�5�2j�2�\Vh6��%Swا��g����J�I?a��������L��	|�_�Q����q�|F) �Mv��j>��6�&):c�v5g���	��e�V��ǤM��S�\[�5E�Z��V���sZ6Z(���==�yO��Z��w�;g9����]g60�J�����J5}�F׳-�Z�=9�-8�2(d*q.�8$�`_�ZH3 � �ܺ��l�������Xܥ��R(M�@��܉!Ie��Y;�E�%�Ԙ����H`T;�yM��ͳ��a�N	��o	��F�a��X��K� �[��et���BW��F���]�$�VK	�Ӕ�Yn��\�Fg�������Vwg���ȫ�]h� ���P}0�����Q���Z�쩷�z�3�/�&����bߍ�R֢;d��+���A���^^H���o�X���"�Hd�#�fo�*UK���?�;7��t�[h���8U^]��z��.�5�sv�����ϱ�^��L~��NY9��{�mD��ZOS�3<�p���������1~�Yw8�E��f�X�.�B�#�!�̭p��2�:9����BR�.���Ɨ�	������^!o�
��-�Aޱ�*� �uu�f�=�
��$+��D@��|3�fe(���8��I�N4� ����R"�H"WJ�)������х&���rUG	�":����`V���8#l�t�J q���̶���m�(t� x���`3��}�������_��|#��Ҥ�����O`�J�]*�j���t?K�]��_�t	<<�a�����*G���>������0:R�"����c[��zn�94�2?�1���V�_�ZE&4#���xi^�&�ő�o����xs��8~���� J��=Q-�FV�ԝ_�)�����Z�Ns|�=�����g�*C��;� �� �����M8�I�8�$�x�ќߏ)����c|�J�Ы:�~�%w�'�:�5��w�`��$UL2�2Ņ2TH7F(��h�C��:^A��|����x��-xN���?p�su���:�z&$R�o���Ӽ�Yŵ�E�v2#B,|��\�3߰�%d�K�bU�_7̀%HP&���hr�G�,B6����d���>N��2��~�DDb7h/D4�����A-��0H�v�t�=O� �P���L٥waf2%��b�A�[I�&6����	���1T��mk��ٵ��"G��v[�Nr0f���@ˎ��u;v��By���� w�MLC)��$_���ܯyHB ��w�1{M%Q黱b�=_*@�5����^:-^�C�9 :�U]��y�@KUyqP߁n#�U�f*}����4�B������F�V���	RK�䲴���j�hUH�U��>��w���"�d-R���Y�y�o0��gw{��^&G��R�|6�L�e��<���.�ǩU���mA�a��A���G���t�:UKv���j:~�j\T%;�C�?��d�$� M; W	K$����J�U���Hgʠ�����]L�k�ԃ��FY��zSצ%�|N�m�̓M>�ݹ�ɛ��w(�o��"ߛ{������6��m:�p{��69�'���N���Y�6�{q5ÔA�)�:�Q��i���j�O�26d_W�&0K�i�q��~��Gg1G"��[/�p�w#���;����zl�R�}��>�l��̎5Ǳ�.r& |�ݪmM˳�g�㳀�u���kr,˱+��}���а���V/RE6�9���ч�ͥ�4�=�/���C�`@a�!`E7^�M���ĺ���F������ݨ(EE*�QFH�M)�+Q����*. �0�<���B�3��U�������>o7z~�����<"SQU ,賟��2��� (���`~�|�k�m؉9��[�$p��)���)�1�$Mo�g�eWY-�9;�0uh��t��8�J�����s�ǻVg: @��Y���͍�O_�Vt�>A��4��H��=�c�u�g��B�@��|]z��^+$\��B�����M �_�ȓn����`eK���_�K�G���%ȭ�ؗ	Jä�UE��t�(E���ʳaqǨ�ǉ��*Y��z��i	Je�9�E8�����
F��z!��i)�i�F���:�P�_�՚cν8F2X�U���袶�7�c����8��0̜8�n_�NoK@0m�Ĭ�aD'�M�bR���'"�)�7�yhZ�Lh"nͯa��5ƺ��e�I��-vM�A��T��զzEoY�XnH���_���X��*���d�Ǌ�V��g��F�r����N��W��0�H�ˑ����gAJ��	=�I�y��&|y����4=�KqD����	:{�����(-��?% W_q�a��/���o���¦	^jIº��Ԭ4�A������X
k26����'L?�o͏X�~��L���!���5V�c����ѵ��Yw���mi$T���C���q;����_G'��u�@c}�e~����S~��|iޖ�(�Q��w;\ཊ�ϡ6?�ȶ�K�ti�K�p�X}���u2=@*�>n�����z��8q�a��zFpi-�,1	*Z12����m(������&�/�Ls�7&~#r<�x�N����}�Q�]ɭ@�(��k�j?J=�v^�[�,�h3ܿ�w�Ŝ4kMU����O�I
>�����6���T&U�\&P5J��W ����[ћ���\� �3�ց�/�gxh?O�!_�B�1㳈_y�}��@"�X!Bf� �q�<���o򝉊>�+��m�"M�� z�Bq�}�wz��9��)����̳)MP�$�e���ʳT��(֨y�Z�\�5P�+����\���)���gsS��8�Q���v@�+�:5��wn�@�O��/F"������&^��Ek��nl
ck�D���i9/�j$���
�9iq��K:*j�^���S�D�\�.q�r��>5a$���Ⴞ��3�L�<
�7���Җǚa��"3?M��K��U�PH��E�����LpԧR�L����l�Eg�����ޏ�ł�ߟ�R�4Is&-�ߛTҳ	-OU��{�.佤�󐹹w��	�ylXx[Y��9
��N��~^.Az:�W,z��'&�K���HI�)T������
 �f-�^�{T���'����]�e�j�^@p�3/�P)f<<����u�[LgϡXr�G�:�Y��b@��{kn7ΰ+1K\"څyC�`A�"�4t���i��LsÙF�0 �����y�vv�i�+��/(�LL'~�@ni�H���,f�ea��ˢ�l#N�ƚY�O�����@�S�p�ėԒ]g�-�\��^�(�;�_'���|��Ka���3��`�����%廙Zb(��N�ʵ��:m_��`��W<��a��f�.��c���N-	�^��C�N���f���p1ǐ3� ��ǳ�ON��E�F/Ey�@5�Y[R��؆�A��}�Q������-�R����~u�4K��f�G�?���݄i^nWBJ��oU��C
���DW�p���/Ups�૒���Ny���Q�L��`_ ���c�B��7���n*.0�ⳗ���+���w'3�{�����8��u��	v�ʚ{�(���h�BNOY�M3���oKr~X������׳}�u���0�/:�r�]��&Q�U��Y��H��(�s�L8��Ŕ���r��N�Bbq8k�8,s�h�+oJ*��S�9�u��1;1�ua����Bo�ۍK��n�� ��z���D�1�6�kњ�	�`klg�F�7�5��d�<2G�N%�ŋ+�ly)�Ȗ�olOl怿�W������>����rv&~���kl�ۢ��m�Z���� �fnR��~i\�����A��"O�AhGձ&��6�άJ��;V�y�'9>��K?I��M)��aaJT�T1MJ��Y�d�HN*�-��V���e��UZ�"�Z�XE[��>�ϊ⪵?�
��E�t��$B��Q�O��KŒug��p�S=���?�02y��2��gd�]����:<=�aʓ�hR}��Il�I�����L����J�u5��I���~C�%D��3�v�KЗ�P��Vc�kMò�r���aμ3T�QN�0�Vm��4�<h'iU��:���~32�Vk�#�cn\�&l�]w�	�X�N6E�� ����VByS�2.XTCq*��x����2�G��*"�Q1
�H�9��٘���%��>�I�
���>����ݼ&ļ�"E�s�_�����\ܚB��	�����lK����w�Q��nOj�5i��q�t�w/��~���U|1l��2���S��jy�2a���OILts��J5��v��Ap�e芝����y�2��?h�t]o�R
������&pJ��L-VN:�����.�ފj� V)-y��nۤ� <���!gE��2�Ș?��K�H=�9�9���gp ��'W��u2Y����[*#J�#�O~'��s&#�si�)}*���iH<:h1+�� ���$�@>��n�\�{ϔ���n="���H°%�^�|�9��&�<۞��AZp�*�Aq����t
�u2��V��L�m�t�q�[?V�<��@����֚gH|o���0R;��?����
�X��O\l{�}�\<�lO��)��dO������R҃=F"cp�$��k>5�?z�%�=�yl��4���}}����ܨ����mh�$h�z8���'�73
�@S96����-c�D/n΢�q��uK�2:�J�o��M�"$��j'��`��Y[�G�����j��r1F�X�v��p�(����-��J��������[˕�vH�e��>�w5�-v}�E�r�G`[x=�|�\`�d�J{G��i��;��R.���fA�+�v�R�<�W�ڬD�fX0�M�3�䶺Y�!�lg2�Va�L��b�gf`�֧j֞���IQ���D(�O{�D�K\m�N���鬽�ܺ*0��M�W*4)���*FYح����������jv4[��UDbE�:����;��(E���~	\�*>+˹x�5�X�D4�}0������Ƿ>H�8�4\����k6��VG��G7�����m���H��m氍�N������4��Q��)�o��0�j&��:�aN�
�� �X ��ӂ�[����!�)"��@V(���6��( ����tҺ_[�Z[�ZSc_�ם(G?(��Ԡ7-�F(�pw`˥Ō,�-F�����Nf�06����y�v#{�zPf��� K^f"�f㰨���UT��Ӷ끬� �u�y�ۿ8>�2_�nr���,}����g�K��UΚ�� �
-F(���|Kl����V��l��� L)�a�u>��@qc��͝"pJ�׀d�u=�k���(�<Ń�h�U�Z<[Z�ۢ'?K܆Ī���m:qAϪ5��<.Mo�~�2���E�ʾ]� �쥻$�H�n R[�B؜\��o*Dn& Y�)��$S�{>L#���@�ߓ�#Lre���􈆂�@��BאָL^�X�L�~է�$���{m�C���p����^s����h����cT���\��Z{�8�[VB����ש������V3�E`[�8fR�+�C��)4�_���CY�|�3�W ������^L��gU2���d���̹ܚ�v�*V��3>�KX�}:����Ȕ�6D! Ob�[GY6%i�g�����w��$��I�CrNr2�G{�hʔ�x�H�z����(VIa���Cl�/�Ejth��U�
1��s.�X���f�o� �X���4obH��V��h)w��g��P�y_bsjzs�n�|����r�r��\�>�R�5_�Ԣ���dZ�_����y�#V�R�Z)���25^�$4	9�nh������MP�G#~�݋�^�RR� s��fz��Ӧ	���c
<;����]�q}�V�n�-��S�,a��̬}�J�H�K-���N&�� �l��ޖ��5[ŀ�h�:]i��#�D����٘��y8����4����v�"z2���.��Z�2�c��}�a��Yc�n��xϽL����`���+$Kz�̽�>�>������IE�tl�54�����>/��_ʚ��x��~:]��pr�O�X��C�*��y�f������A��Y�߆FЌ�d�Jܶ����J� ��*�lE[���,���Oqp��Ɉ\=��h��� ��:KtU�r���+ �!=���m� �#qq�)ۭ�������u�5�6���'����n���yZ�ɏ&A��H�~�� HE�~Ƙ �\�F,�?����?Q;ɞ�����+3����#y�)&5�	h#h&�0j̗)*h�L�c}��o���u����F�[s�_C�W���ˤ*O����N��?�����wԬy�!�iQ�K�����Bt��O~���eA�K�C+�/�!���p5����p��y4�/�	�"�T�b|��Zl�ϻ�^ߗ'��`�b�t�>I���
�A'$�[��4�[7	z/CH�s�|�Z�'��)�����:������\⑫wA�U�'��{�=�k�	���ܿ��f����n�`�-V����̋�-᩾����?1&��r�_�#j���v�t��E�15�p��lP��4UO�ހt�E�#�}X��CXG��0Y{E�k��5cJ���ͼ�1�cs�RB�CiQ��̧_2���GP�W�-	�u����l���F��
s��������S�`WmDWx2)S�C�Y�-�bx��$D�F�;	»�a7N� ����b����"�O*���0$s �
eS�l��؋z���#�q9
g
�U7����$��<qT�߾.��1:��J���V�W�k���r5���m��a& 1%�t�_+�I�=f�X*��hw�������n0�=��H��;�xi���$�1 (�+J<��R-�>az}��nWy�l��0	DI�����P��"�wHń��.�b�`Z�ܔ>i�#ǂb�/�~��HD�N���Ho�/�^X{gSrF'�5�
'���ߙV����f�N��A��"#;�,�����F�	��j٦�˝X*w���;��W<ߐ�U8@�Ej�+^4�ζ��L����J�m@�T	 ]3�
h�΃;��V��_�8v
�6i_IZ�������o�q}�@�5������Tm/�
\��t�j��_��5�˘X�]��j��P�mR�	1���]�����Q�9d�l����*�Z'���H�������Tm�x�M�ѓ����ͥg�t�{����ݲNb�M�+��ݣ�y���0i/����U
�yDr�1*o�r��wO	��s�1g���~�Ex�4���^ɫ��������W���#�OxԌ���tp��lh��a��N�/�(�MymmC��g�d�l��	/K �`����E�Ӷ�!K�ꬊ�ſ'n7SEQ!Y�z��T��s�ˎ�m��H 0���/5Gg��l�E�'��!�F���)��u���\����|O	o�ԙ���B��X�I �'#����,�ī�k��H�ע�b�,ߴ�4I�Fw��J�.hf���7�7�&?rLT.��V(QÉO�'��w�a��ɔ����i�5hP-���N5��S�	�\�G��-�q�^�nQ�������Q�'шn�t��[��v�I�V#_(��c��L�B{ d�g�]��Z�SF��}�t����a�@����q;nC�����#��[�?V:�m\�}*ܬӱCs��J�� R��܀�Sk�q��^$����Ų��~>Vը��(��C�7}DJ_b��u'EL&P�������P�ߊ�؆���di��o����<��2��h�wG�6�!�waK��{��/������&pbQ�e�I���Pޓ.m��C�Ŗ�_��.ZCq�藺Cy���g">�&s����b���$�������I�1ke��!�(��x�Җ�L1���sx���#�ۚ���Z�FG�&������rDi���v>�T㔛��M�ּ��uH��������qs���mC��H���&.�F�^��'n�.*�b�!����{��r�3˜�V�4ĸ�f���|��Bʰ�q��������$�l�oI�&x��b���8t�N� ��a�!�~��p����-	�k������q`Q����YnK�Lz��f���$�βܙ3���xm\���f}��_r�$v���6�#j{>���d��s%�X652S������s�����Ǌx_��)�B�@@%їV� ^b��jN 3��>&tϥ����Su�XPd �a`!�<�O��ͯ1RR���Ձ�K Bhy�T��P�J}a��@�J |�f���b�<E>x���-���sqĎ2�c;����OD���2�����*�W�Hxf*�P!������9#7jk���gȃy38��ai������,�{ټ�FC.:s�m?�=mr8�ߢ�h���I�q�/�1��i3�R�K�Q���K��i�M5<)���>ŋ�8ݎO�e߈��&�Q�~��7ئu6R�w��%����㾇	f�4�Ʋ��*>\&��$oE=�(���nV'�/�B��s�a��ˋ��XIw%.UC;�1�c@�M���}� ���Nnn�w���y���8������Z�QN�,
�t��|�ְ��8��� ���"7G%���EZ"Iu���>�َS �ޜ��v�$c�� �ᮺ��%����}�qR�UjL�|��;%7�N��8�I�#��Xz�r����@������y��v��j��h�֯j�?@9��s��k���=�{D��'��M��SŮ����K�,SI[�[�Y���|m�R�.6�-��2�ׅ:���SA] ���$���?+��D#9ZF���,��oJeϴԳ�����x��#�t(��Ч�ʍDf�T�NX5L,LM��r��.N]$���ug�7�ɿ��e���ʦ�����<��Ւ�m��x�����x���f��<��Fit��h&���=��6�~>���
�b@�[��`����d�x���7K��JP��S��鿱"�B�����é�#��C�3�t�E�n떔$]���0�k����t��eP�N��'�Ǹ�M6���C����_>	�ǐ����	@+�lo-^>��h���C��[3�o��Y��v�������D�����PfEjMo��}�;^�f"w�[�4��B0[�K*�����)�ߗ
L�#>J��^nU��w���Z�2���)�i�FmF�)$�>�~`T����O&��hur	����؜C��p�Hg���9�э���&��@�A�n��S�h�Sc@�i�KQ#�%Dd~�Y� h��\Qo�6��{"�����������?�����R�v#):���7	VT|n�+�x�i��5;>2Ģ��8!�x�H
A��!m��&���tˎVg��
�� FH��>�T9Q�U�<��q���2�`kQ����`n�?d�uG�7�����W�?>�^^m��ѓe���i��@)nq�%�-�D��
K2Uv�q���wk�_���D�Ca�r#~��^��g4��r�r
]�lJg���M���&M�L��2*��;�u�e��}��ʯ���+bc��M/0q۲��cO3�<�v��H�ك�S~)��l�z<����}�"9}��:����[�l\D1A�ޕ�ގ,L�JB8�<����E��/�ٔ���E��x���#,ȩk�Ac=���l�or%q��a�W�Wd��>����ɤj�Q�ۀ>ޔ��h;Q��G���K���kL0�2�\F��z/;��ޕ(�/��ש?�p��q,>5D���D���S.��uF��;�t1́���V�2�c��7p��͚����E24Vٿu��G]��s1\W����{�v�q?��4ιc�B��a���/�UF���So`�6���F|���r�;�8��V&���C��{xp���c���%m�C�KLBn����ep@ }����N�l�2�E�j;h�:��r�D���t%�`����.^VSu]s��B������<΂s�T���!���K��1��C�8c{����b�]|PY|Q/my��Rmuo��CC0��Ҹ""k�L��vL(=`7L���Q�-��(|�wV�Δ�]��l&;�����#�b�L5�XCy��kH� u�|����5��1�W
F�m���p�萔#z����;�]taǣ�� ޻ƪ�H�Ř����@4��C"��K��%)%] Lv���콎��u�6�NRK�@ �o�d_P$JP�9�QA\J�y��\���]ZY�C�u��"Vdbq��V�IN�i�f^�Z�*r��O[v�D���V�5��t���8C�5�:t�I��A���p�i҉2���X��[/��2vǪJ\�[��2���g�~o;֡ |�X���9�162MU��7z�)5A��g�=7�i���fω�A�H�[�>�qy�!(���+�+I�i[m
���{���-��P�>B2�o_~��et��_�p2��O�p"�>��J�>���y���I��Z����QQ���Sx��5��Z3���R0$	�q%�W��k{l��X��2�Q�4q �4>h�#q���At"�'�����Ĵ�dt����~^�Ϧ�e�d9�i�-tvhU����-��:�H<d@���/mz�&�H��hQwZK�,<N{�o�]�I�A�yn� &���_�iOގ�q�)���F�Z�O�$oJ�A�����z{4�N���ұHT��=2��;�s��bCtM����alr0���0��6��}r�ςm���k�}ju[����Wu	UZ�ݹI��ψ��u_��*3V�����o�[pfw��W��"��f�XUD\�j������o�#ErԄ���/�Q{,E֛LTM�+��%��1��� ��l���i�l���i��sy�Xl����z�.�|��rl��7p*��N	�q~=t�m!��t�l/(�d��Y���&�}��s����?^b�0�,�k��$�2�t�l�;k��2���Ɲ�7,6n2P�Szc݇쮃����<^�&�݆/�̹>5�b��$���1C�u�z�,
ݴ9[��Y���m�lк��Y88D�,���,��	���r�����لW�d�����#����wO�c���q���<;
�s�9���BI�G��D[BϠ��H����r��ш�v�n�8�*�.�M�Jm���Z!7��-�F\-ER�YI,=-�bc�6��=�{�^�;s!oE�����J(+��J`Ez��R�����+��ĉkbL�x5��*���7�,�g����7�\�v�|���Q�)�G�G�W�~'��9�g�4M�����5�j�6�f]NNo��48@��. �+e֠�v,0��TQZ�(!'N�ٯ�:�l�f��
jwm�Ǚ����e���>�6U����#���y4 ���_h?��ݛ&���hl\}`�iSѾ���|�N��a��l_o#w����o�م�F�LtV�u.�{�9�H~]�_#�#;	�����Nz��t�T�'��ķ��i�)wy��jc	���h�*��6_GC0lm���Y��LW�0A���kIF�-&�=�l�γ��,��K�n�B /5��bYP�]Eݜy��E�:����ߩ
����]��9�X�.�7�	OO�����<�E�1y��U�z�/mU�R�A����B�Z�.&P�G-�-����fbLE��:�9�vh�k`� s?����ృ���[��"�{^�@�=y�������hT��è|�\��I�M��7˜P_�Q��g2k�a��M}�PR�2�Q�!v��� �.擎`�`��Sீ�Zz4�Ҭ�axTD,C]�!�����b�2�堹N�����r���<���I.
C�mD5lbz��^2ժ�Z��Zoы�h��?�"��&L��!�����ጏ4���qSUh��g�|xY*P^� Rc���X��)����QE�x��u��˗'��Ƿ-�N�����y�� LS�������͆�p
�A�#�3s��V�,��~ ��n\<5�Ǻ9y��=D9�9�.[��t� �k5\r��ӀrE�Y�	4%O�\k?���<G>�5g@��2���Ͻ���v�B���&�j����	�iY��a�ҽ[�?������&��f{�����U�Q�^^J"D���M���o�����gZjTr�E,�Bv3�L�������ՙ�l���8R���v�=�#E�E}�6���겻qt���Z��o<v_ȼ�*t7m���V�%�8X�D3~�A	<�F���+a8�/���F$��%�~N��Aܑ_u~Xm�]G�95(x�mha�(�\sw��
�}\ �6a�ď�CɎ�-���g��^	�h��o��Z7
J"��ST��'�Ӕ}|���O���2{�e���ƦG��v��9(�t$c��.V��'���Dpc��1��d1Z6"��nDH��6)I�����	(f�픛9�牎sq�<=��|b�Ξ�ݱH_[a��(C�������/�u�E�k��k�d��nr=�>�X��r:"Wq�d�}`�@k%��0j��eЫ� ��l�/g�c
���SB`���H�j�����~Y��C�/U��=�	��c�[���$�^�DX���䢋 �LU*�m�\�ڃ	VzCÚ�c�X�4�v�|�ť�S����i���s���I�|�m��Pnӛ��P^6-�p��8=�=T��ǲ�Uu��V �{g����`V�|�x�Sg*�1$�=\�.e�ج�0=������A�2��N9�R0�"S�p@_���s�	<un�2CR�F4��ϒ��&���ą�n������[̂33 )�v�5v�ŊڋB�=�Pa9o��sFG��'��?W���}l���kc]��!��^�KՌ:B��V��#�b��E�Z��"wi�yI$���b������|� �ߤ#���3��'7(VQ��5�9d�M^���8yfv��Ql���gwR_����fI���[�R��b��$��%�B%:��Gjz�vrx9A�:"Xq�D�V�=�M��bY�J�Y���v���ԉ��I���I�#1kKz-���鿣@���d4}f� چM���Ͽ }������B2�F۾UZ4�\����%�bV�oU�	a2�<Ҷ��22���`Ct��V�v��Qs��:�A���\��6ܽI�
��<�f��Sb�#u��9>u\kj֘u��'�W���@�4�pdJV9�f��w-����P�8��t�w����,��߿�"FZh���ʥ�}$�{th@������B�Ib�:Vk�;wX��3�ϡߛtD��ki��@_P��g�q���ؕ��ʩ(�7O=��Oj@�� �1�+DN-�+�p۰���ǎ�x_:�����u
â����a��N�I	��sbb| 3p��A=�)+,�C��s�ιr�D��R�j��Tm�H5�+�ΧmT_�I-,VZSt��!
��q +���1��q������f�*�Kj
�_�"�\z)��W�}kF����9��&�U��㿥���,74]��ύ���IE$����00�m ەXn�!�2i}N��G
5�?ƙ���Y�ŖlH2|�%�)Eo��� &�|h&k)7^{g)��,��8���=l���z/3{l
�G��~L�!G�9��U���vN����Wl��?� �V��N!�hsy�z���J
	r�4.o�*�%j̻2ؒ�X��_��HF�X7�҅�b�]�-Q^5l?%�}d�^�ޖ��f�"�'�ׇy�Ⱥ�i��c�)����(\��=jCjn$�������_�� <P�����
C��W%Y�B�>����H2!�}�P��\��L�xf���	�RTbx]�f&�!�>��Z�� ��Xk���o�}�n�!*��%�ۺ@�fF4ב������*�ڊ]�x��pk��bվ�ck������öj��҆]�^��G��WZ?���/��`��yL�$��ح] Պ\%�w��� �d�I�	��>J�hs�*�	����+��x�a��V(�|;FQ94t�G�+c�ԃS�?DN��r2c�74��Kzy7Hn4R��x�7W��4�.TC�1*�l��'�CC�OQe n������̷u���8�������V����X�����S/ik=E�g�Y[8ِo
ш��-泶�e~����9Jݭ�X[�O�7B�2H���N"�~mY:V�`g;܈�t�� �S��,����,R`s��U1��bZ�%��:Tw� �v&M8���U�7����/66���Z6�/O��C�.���߽�����[ �8�K�l=���Qh�!3Ay|R�!R>�<M�֋l�
�`F��L��z�.�Ҕൺ�LD��5��9�u}�yY��D��^\v܀3K{@��̾��I��*����!���{Ư�1��r����Or�	+K����ɸ�D�����5S�xn�)�JIq�A���Y��W����m'9�?�'_c��Ůb̷2��k�Z�����������8t���~���{�m��������XU�ԉ[��(����%��)�s|����q�һ&�%�~�����>�%@3Q"�nyqC��#�eW�?��ZM9eُ�����wY	m����ߧbu<��,L$�Z:�'���h��$���ѧ{��B�=IȘޤRn"0�D��H���)���4^Ѝ�Z�Ɖ��c�s��S�@�}� f�%
�*���fHr-Iw�m0�!��8��SS@�O����+v��V�AA�/�O���K��Z�k��u�����}�˧�J�ai|ɰ*��5t;bz��R��U%ٰ�0G�~&� Ų$!��L�(��c�wߌ�.�e��R� HL���|6�+���T�l=��.9Z���T%�4,�O���P~A��S���f�Y��澕BF�!�����Շ�ӄ�;O�S�E��ܻ<Ҭ��4��af�Pa�Y��"
O�V�s��d�콥N��&�|9pX��X�����) !'�1z��h�O�N�Z��� ��2?}�F���d�ښs��n�����"kjs�ܽ�2fU[�3�vpJ�J���WD؝�*p�S���e��5�ˑܧ�� ���3)�P)Z�*v�@YvH��@{��qˮ��DO,r@1���R�v�6��2�69h�"c�<_(�	*>Pү1'E�I�7	�}!�^�	А�-p�� �`�[-|�p�n�̷�P�W�!��3�ƏkD��A���9�a��2GJ3Y��*Ԃ���ʲ��ӛ������S1PP�$���b�/��:��&M��Ú�̝�0=.�
9^�V��;�Kی����揺�4���g���kv��� �$�9�t���6P�b@N��\���g�P�"�g�r�u$y%��Z�-�o,%{!��iω��lҭ�&�	��?5���K7*s[���H]1������K�?`�����,���[_��׵�s�C]�՝c�jZ�ľ]v����ۅ�s����lQ:ù\�D�w��r�K��=zHω�jyo$�Hg�䵉GW�D������E�6m�Q%�뷦�?Ky�_/k�`�%ڑ����)�6��r��:`�U�����nK�k"�g+�5����s�n��Ӣ�^l��)ø���(�\X�#0�"Qy`��_�f�d��3!h����Y�6E�v�!K�0@�s�<��٩r=�0lN֨����sK��}�`2!�Пx#�O�z8�c�oo*,9��X�A�N��� 12n��}X7����3Yzf1�IG/nfs>����"�6���d"-�U�R�Q���ʬ���O�v^��"���]s�����SA�B�t�{l
tkbC�ES��Rs��vb��y����
/�� yK�?�>=���*F���K��1�q�;��j�����C�X�w�[��y�"�:�O��AU��_�Bv�K�G~6�5Ud��H��8Q�?�<�N 6н�e�5�p.!�ٞ� JP��R&3'͌ ���S/C����d���\��	MQ�{��t�j�X8��
��kE�6�w��֊Y����<�8�0[�m�,��R�<���@=|��2�-�����|7��Ԇ#g�|�\�4�eeR��L���%~oqٲ?���&K�R9���&܂dŁ6Y�c�x��ղ�5� yL���`L��~Vՠڵ��S@7��7����kfW;U�B�&�ߴ$@4n�KU�E��l6��Բ�-^����%m�	^�[�����Т���s���aک�>�[�p�r�A��d�b����j�* a��1v~νk�k��1��5�B92�T7�����5o��!6
q�����Pd�_��u�2P�=���A�ag�~���h9:�@���H�1/
����MG%�����c��(�xq�6'HT�ʑ�?�,R|q�B �Ms���5Y�-�4����mz�5�?��:��;��S{����W��P��Cxy_�p�@�^0f����eǏ󘖉���Go��M�v(��o!��!5�$�^j��T>S������}�����U�����.9=����̼��)Ip�N�2#.� qM�j;�6D�߉�s��/�����w���= �ό�+�,���؄�bR��l��ņd�L����˫����/8D �2�F1��1u9�p�dz w��o�Mc�k��n�d�e�����"ܺ�e;e�V�G�����s�xF��9%UP���ja��֊�07��_�<�ɼd�x�Oda𹢕�l���F4%��8��Q%��S�D:�-K�h<���OMP�x/���s�Rؑ�;<B�)�n)��#D���նhj����k���9�d��`~F�N3���f���2����>K�T����=�3�����ڬL,��0�a#4U���A�O�(�2I��LV�J�R���<�6�T�r��k�Q���X#:x����H�(��RmaPYkJ���t���^��Vݐ���'_��c|��uɅ	�^z���IʵjlɌ�y�~wq���Y���0�����S$��<�KS!	6P�/a�������p�"܂���"d�Y
�=G��h"9�Su�ח��\!O��B-,rUNn�ߠ�U������
G]��O���ȗx�������qÂ�������P��:�/�:�d<`�<�k�y��[#�;�o�G��r_O�>���i�������ݨ�nܔ3�-������/o ���p�3 �@JC�!�W���>�!���.uA8I�k�GJ}7�Ő�O8J,��$:��uB6�eG �$R����{0ͭ�E�"��E*Ns1�0�/�fw�`�'WM(P}tY���NF)nj8�E��$�g�*��g*t����L=���*���	U��>!���à��Z���3�3�f	�J�@U��f3�0/�^k,�6�6�V�����M#^D�۰�"m{*~@��A��'����$:Yw�#Q8���@
i�&#ήg;F�n\�W"� py�W1=z�\N'�B�No0�ĳ٨_�'h[�2�)$I�F�mMl:ӏ����J�0�E���p���&~=�Uf�30Ǌ�D�G���4���vu���f8i@�(��D�B�����iB��U	��4��ɒ˗��\�k)��qo��3�������42v��OL]���#T%7_�Mm+d�"���2�CE��:�L��Z�X�#<U��V��pȇ��k⟏�g�KSJl�RX����M���z:�+�I}��xA�f��H���<�l*��ޤ���N����ii
�?f�ӡ��L�2!�H��}=�KV:.���(���`o����+��٫7��Z��W��<avU	�ê-�O4��
�d.
��/zl�Ȭ��_�7 `�U�|�^�A1 lV$�.nh��6�;h'�d���!z�@���dq����?���[��s���ԓP�E�.�(�;W��:D��.=��}q��=NE<�)��5ʏ�
 mp��0��9G�����dh?7�\�{{|����P���������I��;%�7O�7��XƐ�Q#��]0�Н���23�}Ħ\&��l��n�n"��|�ϔ����j�Ϡ풬�����1�pZ9`�ܮ&j��(�)!V��5�y4����y��QW?ɝ4ʹ��*-�N�����d���܀�[uZ��AS���HW��h:�T�?
 ��d���m���q�==t�0�[<�N���2 ηcB��� X)ҙ@��H�k�l4Is d���PYu�2�|.D��m��ԭ���--%I?>{�>��A�@r�z���֊�񡙠����A�ma�6��'�r�� �����U��h��7�KL�D��+:���"-�L��6�l���ۆ恈�H�O���j�E�߰����[s�2��������,�I�����gՁ,�^��K�+mÔ4c)�*�z�w�w����d�O6��j����37�ni���}��P��J^=�9�V6�Ҝn#{�!��/��������t..7Jc����e���[�!x��8JB�k6��#�&����@֎��{�4���Ǯ�S_O�ll�q�L/l��
2\.�s���7)��ކ��Hx��n�;R�=��-A��Ve?W�TSPq� bos@U��^('_�տr?yr���Ե/(���t�00٣^����k��Rnsev87
`�C�Cjҧ$?I��|�J.)��Z���v�k����N�������C�dJ�b�徦5�Ŵ����Z�����qgJ�������b\>{q�J�^:���%�G{\!{��@'1 �g�D���jD�L�
���i���X>wP�o�F����笈��w~�V�P�~ox�i	潊N�(�%tI�Uo{W�}�auƍ/{Y֬�,(ss7�%��qZ,{8 }n�n��3����$�!�}	�'���W9��*�bmK�E�)K%��	�d�f��������R�qX/i���H=-|��)�����B-#��� ���І8�*r\�~�PO~��a��@�7I���j�{����Ϫ��Y��\�_gF�Z�g`�]	�9p��Љ�kӫ'�oDA@4`�	=���aJ)l#�7`�A��h�5��e1�w�pɀfн�l������d��a2�� �?{:Yt�C���z�xw mI���[!F�8lDM���z����i]�&t&�K��;�w=""��	S��_#9_u�ċ�4܂#�� �~JD����7φ�8hDs��%�^�픀�	P�;!�6�CkPztFU��L7�m],*IF�S����+��^œ6�4� ��'j?S��`�S�+�0Ke���
����SN�ݦ��Me��x�mڕ&t�E�5>C�*`�=�"�K����$z�M����iQCX� i�#��~�������"��g=��L��K���6�Vy���:��2A�3�|�"��4kh��(#��i�h�sC4��Y����n.e}�g,)�J�q$:�;�!T+A	�z�c�*�hq������C�/�����zOXp��_�����V CȌ��V#*ر޴��]�7KN�����܀dK_��\jU�m��c.[��|�� ���.�["7�QMа����)���(P��>Cz�Ws�z�2�7Ы�? ����/ ��o���g>��8�Y��V�5$��l�U`�7a�vvz ��7�|c4�xš�o�,#�˛#�LF?A��:Ƨ>�ySm�H��=!�1�@�Wo�S�l<{��b1��3��΁��mD�w��F���KDj�h "?ȝ��:��S�6$u�5晌���L�Z���#��yVU��qy���#�E�Gվ��o�ͭ�����{���vF�rO��m�V�<���4�#�=Fe�kS�m ����!�`���^+��A�뫿��X�.�NӨ������\�=umEaO��{�WW���F�U��1{i�}�,R3h�2��<���q��y\tǱ��D`{�����r��r�����q�A���a��i�)zj_O��'��Uh@<��������G-�6���̍|��hy|Ѽi-V���r��@����:�3���B�;�=��0�����~�g�}\��TdYj��Xࣘ��&��fizP�W,�
��y�4~�5�%�١qN�������q�n����#Р��i�7-$\�B�(b�a�8���X��^G����ɆVf�6���a���[?ج�D���B�fO~�<���<�<�A�57��<ad�������3����dy�R��a-4i FKcNo:s�^<��V�7��j��1�1h�PK�3nG��1E���4T��ip����X�x1�h��/8
�neI����Q���WZd��[��J��z�h�2��t�p��`��@�܍m�ޟ���zG����uMBx=$N�F�8�8	Ic�j`u	=�n��9�i�{7�8�}m���d&x�
�AN
��� ��O_@���x�5K�K.�<:j������ ^����12�68�oZ��ASy7�뻚� 	�nF��9�"́�l ���0���T:ؘ�Y�5|�ݾ��k8���m�s��8�NǿT�S�2ߏN[_u1�-t$�'�o�hh��''P��L�9wS��ʴi����PXgle��m8Z��fS�
�N0N�H)~"�)rM�um���5��rޑ�b�*�M����`���9=<w�s ��g�ƙ]M������<?���Fs!Q�$O�Ǳ�x(�L������؁Qg�GT��u>�X�~Y2b���S���|)��E��R������v�
6����j��
`��O^�u����S�~xDfWQ|����j��@��t~{"���Y!�R%�)�~�(�"WY'�ґ$Z���k�*?T�k�t��4�~� 6�L���j�ߪ %᳿ZHLvt�)m���}�(�=�+幅`ͦ�t}��6t��"�N���䂙��S�~���0y(@g婭qW���p�	dG��J��S�\�k"�2�6'��B��k�&ݦW��>� ��3��1�uv&�e��|C�!/WT|g�3p�����J�c��"F�b�e��R��	�9 �1��ut��"���O(�X�ӮY?���q�79��7 dۆ)��TE;'T_�������������X�f� I{~�l����a�O���޻	o�} ���I��H LI=#vH& �?�W�ٯ���&FO2|9��k����Y���=/�ٹyNy�X��#�܅����:$��'vU�e`�U�G2��"�\�B�E�p��ܛ�x"��v�EG�;§�`�Z�C�~���:g�[�h+��Ď
�6w\������Ywc�������f��pǅi�M�}��m_d4��=�0�w�5��H�#�E�X��:C��A�\��ղ ZP�����IR�X�D#�齨��G' 3#{�5L��=f�sߙ�L0���Gt$�b��ˁZ͘5��x��!�6����"zc.p?Z��W��;�qQ/o�A�BU���2i���8��?!z3�z���q2<��?4��ZZb,c���xF��1�_��a�	P2��`0���y^ы�����ɨ^m�ً�Klf�����ܛ��m�R�TR�Lu���}���h�ۥ�,E_��W9�a�V���d(�Y�b�䮷�X �z�[�c����x2�Q���FF�,n�[�$i.�Z��j�KUa�F
^H6g��n5�HDc��l	j�_O�A�W������?\��39��o��=̑FZ\7��!;0�.'W�%iQ�1�� 0�{�q��������0�_T	eq���F�H��母��̒�����]�!0p��O�R�����N5�
�m"�7^U]C,8C�g���ߥ$�o~?�;�<��H�M*�S�
�jv�4��7�:��g�c�E(�kM Φ% Ih��/]��ʗ������}��V���DL�'�8���V2���?�FQ3�8��&��vd�䥎��Mt �"����g^�Bv�ə0�+O�� \�Bbez]`� MI�a�����·
�j����Z�C򥵲h�\u�IG�2W��<<���m'J��t(��P%�𯏀�3��V����Z�fg�a��V��ႀQ%Ģ��[!�i׸b_��'�IU%%p�u��ե��"�>��T��ͤz?w���Z�I���t�L��2�x*cY�S�g��q�-���2s�C�9�;��og^M8��b_��}c�
�Ǣ+�!iw)=K�(�5z�7�C!yƾ�O�ӏ���Y��9�Y���jil+PwՍ���Ct�
N�/� G�m�KP�Un`��m�Doȯn�鈙Xa��g����t����L�p�q1�.��E�i���"��]���Xt�1#V;H������6�`6��8�,X�g�[S"Q�jUak�����#-�b/�	u�DWK/����שn��o`�DN�?G<A���L��4 �=�|�F!%�wf���l"K�����/�<�k��^"T�`�;e�Ch��JV�x8!�r��D%������x�ȫ���{��U����4���M,�@�u�(6��t.�T�49��Δ��)�\B-���Gѱ҃�	�����)���}�;7qt�� �M��,��\&#�*��zz�@=}��*]��Zs���T��}N��Q�+_�Fn?�@4[��鄸R�I��}���|�<΄g?eEE�R{��e?,�1�,"� >���C�p<5�����-P�Åj�n�b�����O�(���7?����2�Qw=��C�E�.��UG!#&���2��Ha��e뢝�J���\�26�>"L׶&�����D�!�6y�78�T�@��r�j�,�'�X)��F�1�$��Y����T:W�����p�,3E�ޭ<�f!���M���Y��eq(U�S�������ʃ^�Y�]��
/�$���g�~D��bVխĖ���|�^Qgt,Q�LU,�Ά�7hx���"��H��ԛ�q��f�>n�2>r��ͳ��ݗ�!��B
uB���IO�Su���|�2��5_(���a��d�J��GH��w�����1~�!�����1����+o�iL���cio+�+B��Yp�	m?�!'T�]5�8�4���k�J��L,�ZBث�t���f�M8��g�I�a)~�D�Ai?���rR���"4�L-4����	�gXa�v�%�И���i��)�h��5����n�W�E����L{�q���<�k�\x)��L�@J&�
K��	>�.%�����ǜIe���IyyV��J�^��:�@�so�0w�Eb�b$D���lKO�:ö����O �sa_��6�%d�!59���tSxGaֿ-3�j�"f/���cT�@Z������j&'=�7t�n��R�35�	�$�!d�.�-�~��[�m�8�m����mֱ����4�����߶���z�7��;ݗ.<Q�*z�=9Ƥ��Z���G�-@"ބ4+�����A�-.�A�w@�L� �;�I�8�-Ӌ�J� sv�����#�4`�]+����ҳ9 X�^-�}d���uuњ���V�Q[9�uء\�+���I
�:���n�����åN��Ĺ }�zi#0��@d7#���:)m�8-���x����|��������������]ӀPI�^'�7�B��W"HJe����-��:=ٔeӀ���[����=1���ݩ�5��K�AäQx�q������l�T�P;���3����J��*e{�RZy5�qb/ؗi�S'X[,�Q�n�H�ƞk����V���Q��{����:)B�X�3SX�	E�_.��A�'w�x�[fs{�8�{Q�������2-՗ f��v��N�5<f�܁���2M�����E�t�F���2^q�;�*��aF$���6j��=o���b��B1 R��Y������jٿ[@����?KK�ڒ�HnR$4� $�H-kt�t�gS�s��a.榗�s�ipܢ��׸,6��W������m��NO��r����2�����"qݦ�6���{��.p�+�-د'�7�8iKO���2��kD3?�D��3��e4?c�\2��}~M__6��ƑI�ȫ�S�$l\e��ũ��$�#&�D�'� ���hiJW��]ǩo���,p���D+<���n�_!pd�$�X����Ŷؿ���j��f6f	m�[�ٱ�[�zx�"?�H���������M��E�-o��M�q�NN�`S)f�9�WioT� ���3�m:[����Ӿ^���oR�9�����^A�����y��blvF1(4P����K�K����j�A}�
 zQ���JnS�� �.-�2fa_�I����R�Բ��y��ý����8l�H7�_lJ9QA�c�ۀ�֒��یaAQCax��&m�Z�)�������6���ށ�������9��c���J�L���NX�p��߉M[�R�F"\D���$R���=�5����c#�5�>ޒ��l��2.�5�����1�MJ�#�,uk*��[�,���4�J\�5��qsd�0���qsdU"?N�gR�.�vZ����F�2u�kX�9�Bq�ѦU�(��U3@��:m �+q"���-s\�I��z�����j�8�����KK�v��ݞ�����NFoj�ݭ�{%ZH�̨^B�_u\m:�Kߔ,А���x����l���i�F`��q{5�У����[��2͓��$hW�-&����aj�vR��y ����*�<G�;G���_H�Ӳ+���-�6I��m�h	s��/���d�B��c�o�F~�{}L�̽\�t��e��h�C��`�Ml�i�����ܲ��X�&��g�ޖw{�1Kd+0����e��1�S�a��\�j|�����e����&=l�*i�S�(>���nk�/-� ��V~�0+4cXJ���o4��sT�n�cp*9:��������i�"VjR�A�NV�SJ�������O�7/�y�-#3�i�u�B0���TbJw)}�++�sqし�� ��X�����L���qK�k�]p�kv5ᾣ�:	j�%���H�}iI���<tb4���Z���l$osK��o?<Y_��~)N��	�nΉR`1L������r���p;&ն��2N�{��'0fYb���U\�On�}�CkwU`R� ���S��Yy	\jH|%�+ ��t:��W��)��k�!�7B���p���i9��Iǿ��(�MiS���,��0�WT�1��rǴ��uL�+G굼!��Ȝ]$e�b�C������+�꿲�>�ѭ�A0qKl����Q��-�	o�&+m�tOLhu8Lzu��5��|����i����XX�#G���&S9&��5$�T������FL@�O�}��ȏ��9�iP��o\�,n�𝯔{1�
-n2 {�H7�S���c*h<���+?n�j��HĽ�| KXaK�[�T04�.TfiS�l�#Ǚ��`�yj�Ԩ.6[9Ƭ̇�G��	q=!�-�r-<���5NXX��T�D��F�v�v\A�|=��Nh~��V��i�v��V���ڔ%)��ƀ@�VtVG&e7B"���~�Ldvż��7������F��B�҉�{���V�=���J��:yO|c����\Ш�!���Z��L,��o?Noo�&�4�g�����7F~M���B�����#�[��p6u:҃/���#��Z��̷���geJ�<�~���!�mz��GA��*�>��$�:_$}�8˂�q�e�xN��Q�~�kz�۵�E�#�ս��?��5m�	���k,E�X�3���Ms���� "��Q�BzL�ܸU ��0�5G�3ڗ![�yj��?kR�8�+R0opX3K�ǳVp�l_^����{"����5�@�Ρ���.N��W������كھ4��������ZKn��@�^hqaV���)�>G��!�2'�2ٗ;b}Q8�v2��E��NoU=#���L�!��[��`/r�w�Ý�ǊǝU�����AN ,�O�Ǯ�rИ߃uA]pً>)?�*.R���:�IU�`Ƿ�)���D���J��J�"h����F��e,К2T����F�^����ug�&��e}��t�+�<�S�6��p�x�m���V:���KZ��g��{���$�Ԑc��~�L 	��R��Y��BC�'�p��?,۵�G�˘�Ad�[s )��G���8`��l�/�e}:ٱ��2�W�r{�9^��Ժ%4�j�Tv8�m�SW��T~�E�k�����w��/	#!�TM����`l��k���g��s~��� K��|G�yM���(d��K�e��I���=�d#_���v�|��i\.��=Bq���m�pn<�P��p��W�W?��s�67J��q��6���4�e��plra�R��*�@�V?]�6���=�܃֑q�+F���<��
�@���N�_e�h	ᵔK��t�%�e�^6S�'Z}B`�����E.�fu�����kF�?IӊǤ��X�ڦɮ�7o�,�\n���38-�&�PҚ��oOG/��� %���͞#=�k~C&|K���gF�%�m�v�6lI�''!��Ț�lX�ة���gY	@�+{iq9e���"�W����5���j�*Y�]�*-�ׇ���,����?k]�i>_��k��8��?�g�\0Bs�t��-?��OI0�~�W�9�bߧͮ3��yz�1~Z���ץ�U��.�iDh���s`�M�C�3#P: �Q��&�-eȘڭ�|S"CT�|K>qr̥sxf߃�ϊGB\�a�S��f�ztHv��\G��L���R-�?~��,�.秮<����/��]�W� ���ʇ��u�1挵zX���b��0Q䫾��vB^�^�0�s��$}���b�b�G~@�[N[@f�-�>~E�]~�>(4t>�r��5l����V��ρ�	0|Vm{����
��O��O�-���lk&�n�����@���u�y�)�r��k���,ZF�R���3�<xq�(�_ߎഺ҉Q�S%����;������-�@�f�=S`F��"�#��.��[����E��,��>I����!Ѓ7�3g�k�ڬ����lc!��q��&�"�n��&!X�ڄ�Y� �$a�"�����Y�z�PP9�l\�P�i3�/ҧ�)(�F8Kyaw^�\�(���X�E���n���T
;9<
���Z���!R鋒��
(�~]��(����H2k�]@����ւ<�h_�x[5�vVL];��5�z�R���!�w��9�� ⫕���z͚%h)��Ǣg��
*u���s���(@���%�v~ec0�!�L�b# �����v�ƁM	��������)
)p�_hև8�EgQ�^龥{�HD��e����㙞Wfݹ'��VȦ�eܖD������ӫ���Є^����_u���?�r*���6PҖ����G��iaz���R�+p��)ⲳȘ�Ԅ�0���)��������4�#OB��"rL����
�� Ϥ�vT |�����bP�0��x�zW<�ʦ�G4��^\VS��jl)�^XT6.��� - ���wU,_Ǽ(g�.�$�
*����Q��BK=�|�]!�DY��a�4y0��� (oCpHΌPɑ��Q�*&���]�	���E�2�o bHtь��NE������6�����}f���X��ބ/�$x$rH+���'L��J�wF�z�=�a�6ғ�i���Q �����Ѳy�c���(����M��G��OA���?���CpA��=�@Ɓ)�H�r�&��Ϋ7�t�w	�j���x��x(o*��EADnʇ�\���S�H;2�G�2��d$��t��ɺOu�(+Z�DH�ŉ�>�-�Oj��-���������=�w�(Ĩq��;�`����
��F�5yl�sʯO�%�.ER���Q꓿�#p�2��U'�ʻf�G�(��I�I�D.U���v��	��~J���F/;�=kK^Ń} ��6�i�.E����W�/���}2�9H�K"��	��_�Q�GK^#U����f�ߚg�vR��iQ�5 tQ��@�(��ܗsU���),}^�°�e���f���{8U�.UL<�s��;��B$�dw+RT^�i�Q�^����g����-��H�?^�t��S�!�.��f��.[��u͡�{��?��Mb�p5Ĕ�ϝ���F+���Y_�W`�h-��9���O��i��+$��#L���-iӇ>��f�Y�*��}��V@�el(P,1i{�R>' 9K�d^7��8��-�yI0B��&i��6,g\N��5F��9+�ag���%������td�N}��7T���d�WL��JbJ⟫|B�0�p�^7|�l=��N�(�8���ú��6����� �q�GR{1���璐_�.5��Nmoӟ���l^�C^{����	)�ַ�UiC��aF�"0�u����/�)�!ɱ���/j�2�^�C�D�x[5���z�e�<����2��(]q-�%��w�~��NM�T[���v?�rz\���N</q���*�oV���8�M�,���/�[�|}V�n�tE\��J��Te�\_�XER;]J8����K�JS3�ż<��#�}o�m��Sib�8�K�>R��
��/�J�y�!!p�Ƣᱚ'C��TP@��0��KM��Q���V���C��.ԑ�t��j��K��r�$۵��H�����u�ϊ4��tt��cۡ�|O�K���Fƾ���A��+�B#+�X���证h��p>��.KB�ޢ���J�0���JH�>p��e�\*8BV�S͋ʦ��^�_��!ﭵ|3_�}�g��q�� �^��+�,+wv��~��	�G�I�-�m�*��ܜb�F�z1�Y4�1F�G#_�&�)����o�*ֽ���8?��t���r;uZ_W�S�c�����|/|x�N	���n��L�:Ʉq&u|ǉ/����on�%W�������)StY~�a��{kq�I~�J�X�~U��w���,�0α��V�˜��"�b��%�#4���E�y��C7٠��K�u[LBAF�&/�f��99�+U.N��HwX�9�GR./�Č�Y���S���X�ٞ�_Zul��`���(sv-2��ǵ����q���OT�$2��������#0+��]G��U0���(�3i��Tj�f���  ���~��1�I��� �i�,��<P7a�=���(RΔ)y�9ʩE�,"�Z�}��M�,��}��/e��hF&&���7P"��J��:��w�T�=q������[��A'XV��F�6\�W#��oj�;[X�L�x���V��0����<!�}s8%ݮ�KLӍ�Q2q]C���I]'^�8��u7p��v�H��=0z��w�%��fnw��g���'�7T��i��o����wg[�q���f8v�+�A�[w���L��0�Pq�E�0�z���Tj|�*��p����C�~�vj��o����&�9ɂ�km�:��i�@7:4&�%ܴ���]��P����]X��4�j�3�h䗮M�;�ޱC�yr����@^߹����Ղ/)J�2��S������:���ic�p�������B�T�7Z�6�:�$3���ߑ�|P�`�Z��\�O�f����c�%m1�,�*�� >G:7	)�W�H_%�i��oQwd������pMlX)�TY��=�=+�ˏ4��t}����٥|!�o�4��&��g5-o�q��4*������u��p1��DFl"4�Mw�g��:O����k�t�"����mS�vCGL���V�:/�^NP��}p����9J �eOѢ�V>|��$sB q�C"d �S��d;�~Ki�W����	��ƱX��=�
q�0���}��K������"�xcW�T֭d�		b��_�b+�,S|*!����3�� ��aOc�iZW�/:�~�4j�9Cޯ��З�Q� �Y3�����˱\>
Z�C6F��=��g1�Z]s�>��iO(��3�t�����d���=�I�*��5B`WQ݁mk��uO_�̓=�[s�Y�|x*���Ƥz���[Y�&F�:�J��"�]�%� $��ޖ|��������K&) N��5,o�:[Ό�if1�U�'79_�>M�>���R�s���+^fN����w1.U��p�M�.�n�q��B��*�������^�����z�<+�F������@�2�������UL��$�l&��h� P׏4�
�s�D�[���V��b���+���ߨ^�0�6��I_����0%����#*��s�Ӗ�1�cc댁�+�?��B��0ƍ�ʡ�Zi����V�te��@��
��Z�Mˇ���O���Y���+��Z��滂�m	�h���4]�Q_�����N%_�δI["�~��Mn�(��t�1w���$ۦL��1�si�KwJ�*À<ǔ�B̪����J��ko����p �F�<|3�����Q�>ʏ�������3MȤ2�D��Z��ު3~pAflD�mW4��!*���&����/�x��m' ���?,T��p��� �!��|�e�ʓ�+�d<�<�s��uk�;|KF�e�h$y���B��x��Lq��;��(�m�N
{^W�J��;o�Wzl���fy�}}.z�)���{u������U�{~����}\�Q�&{F.Bl�6D��d�cM}H̢��� *�-	�)����[�Qt2��u�N�EcAl�N=�U�F,]uŗ��v�9�a���>�zf~s�e� }O�B0ґu�}�W���j�2���4��s'?7�����3�\��\�����:CqS��ձ"��RѸ����l����X~�-���&����]y��Q�)	�ޮ�7�f��!������@y&R�]MA�䦕'��U^^��v�~8J_�M޾�G��JK�U�i6�N���]�s��$��1�E�W�%�%�j��iח �3Y�����wT~�c�,�E��'�Z��po�"=�l�x�j�G�^�O�L��[h']��i�.�T?��5�� H�E�藢�o�俠b[	`�0�6ʲC
Z��"��{9�E���ܑ�_�ErH��x>�����'mA&�Ѡ���?3���R>F�����1رޱ�-"9��|��f�BFS�)q�tXkuJ�T��"wW=�&q6 B�=o�TxX���[dI�#4v��Ȧ_���lcjܴ�6���ӻ� 
�G=zAK@�{}~��V�5;�^B>���AɾY$�y#�$�ǻ�-K��8��X�P�.���`�.�ݷ�vqC�dK�g���#�� ^;&]e�������$��&j!��vU�C�@ ��pAƝ�2��Dk5h_m�	?���6�T�H�	��w	ݪ����e��ұ�٤�b<2c$��6��g479�̹m+JGҖ�ެ��<w�V�MRo��0	'����O�x���Z�S-	�cl`X~�|���>�pe��f��R�EǼ�3ן������Qt\���,��
�I��m>1Ćxk��2`�nFNP���/�r@P%����͂ Zy�
��|���8�	�I���bn��6���S*�V>[J� W��$t�'��M-��6r��䱗�_ݻ�¥/��$d��O�ZHP��ȍ���HY'�M"��|���Hs/2.\ aWՒ��ݩ�#{s���:���t��)3���7X؏�E�fJ�v���h�h�H�$= ��L�}�O�^�4�A'�Z`�����
0���s,���k<֛T�I�wf,���� �� Z�,�@b��TE�m7����/v�p�m.n�q����ĭ@����c�t����V�7��W'��~'��M���Ee��\���kW��EE�)�~��6���O�Ȑ0S��xhdL�x�.O?���R���y275ʓAZ��V�SOYsdu�D�GG��f>]_W��MȊj$���'
����W�'�ï��S�H�fd���n).���E|)��+*L��SO�B��;F�X:��ϖ����'J��.��n����y����p�R5�S��EƉk���pϐMh�G�-��UG��h���P��o~��u0{/n-���=Y�n�e���	���ٓ��y���ff]N����JX��'�ۡ�}���Ds�w0�;��Z�<i!3���*�m��k,�9bg��ֵ���J����7�^-��R�����)�7D1iHd:�a;"	;]����u-ߓ�	H�.&���Ł'�i1�!|�:2����kH����T�u>L��)�0� �>��`N]U�B��n�edE�uқ���׋�߉;�L��j/t�k�-L�'JyH7�<�����-�W��봷re($��x��Ip�f�?�y�����A)���>���n��B����	`Tmo�7
�b\'*���V�VT�ȩ~=��lm����&O�4���,����R��qu�[d2�.�q�Cr�Y{�!50{�:8�-J�L|��0����b��y����i����30@�4� d�i�>��K�ūC���i;W;��ҝG�ڤI�2�5�~��!�}���&G��ӇJUr�lAF�������� ��n fN�[�v�%Sv�k��l���
腯�} -ݞB�n�7}�%V�a�go�� � 5sc�=�"J��Ļ����'�[$��^�%���A�Ů;��3���l+�%#<cR{�	��E3$� �/�I�bx��5�8 �c)9qQ�6����PcV8A���lxͬ�����\3-�C���Dp_V�v��"��S��3AC�;��E�-�����Ak�Hh|��
]�vw���.SQڇ�F�T�{r����(��)�p9nŀ~�}A����V�����k@����_3��/��L���T�M9�����r�6�r��H7Y�%��Km��Q�
�%(� �j�[�oF���Qa
�ޣAl�0�C����}|W�.[A�9Wpm����f�&�<�|����{T�9�;�S�L+)�B0��Л�GB��J�u��:O-�|�nÿ)�-���w��8����B���W&±'�iÙ���'��$�� �A�������������2�~�swշ��QwK����oK�Ta�A��6�v~ׄ+��E���t$�_lF�kx%Q�mKy�o���ݹ)8���N��L��A�{�Ã�E���5�
p
6U,s��e1�D�>-@�_b��)E�T�
ZA��[Z��Ȟ�F-���vD
ǲ����F�m��'ҾW�����/�LB�C�9!��'b�� �o���-R���IX��?�x�ipl��[���� z�d{F�aȰ0/���ms4���e���uU{�FѷSQ���QD�;b��q��H�"TE��	�)杳�y}p3��4S;����N�b�F�F��w�'�����=\���̐[�g�G#�:��bsd����qGw��a;3��'�v@0�rM��F��M��6���K�Y��Y��%d�������I�v�T������H���WK��
� �� ��J*
b2%=���*����_��&b����)�>�A��d"�0g���#]��!�:n"�d� `�5�'$w����y�wo͍i�(��e����-���ע������
[5�����>Q���RT�֐�,Z��[]���bW]������2?1�	�C���Y��q�b1��e��8'�����Y�K6�`��Q�R骍 ���-�6	�*��h�--"��u��O���o-ia�ar9.|88#X����O�����U<�%غ�YS*�XӘng�L�/2tVw�e��A5�xTN  m��Sc�Mg��� }�J�0��{���|�Wފs���<����]l�6&c��d�/���U����:�����c�e~�9��57��*��L>Z���ES˙tҳ��5=��8_y� �TӘx�iؑm��HB��p��r.
ú,v����>������L�R�������p�Z1��RFj9Yr2�Z�W��6'6d(���U��!�f�,sB򘅺�h�B9����JU���gU[4���!��x~$��$����o��9ts�m��)�j����1N�"2�'DKt��U��
α���H�ᚋ6�[�O���9<�����v!�@�}��?+�]-Nu��QL]��Vw��E)zd"%�E�̴�OsY7��Q��$��b��h=��g<��aօ�ߺt�{ڠ�-l�딁ff\ҩ�^�Qr�l��/-%�����$$Xɶ�+���Z��M���}E���u/��4Nǉ�c\��~�˷DA#��s�w�-��^�~I��O@$26U��Y]��/>u31�j�.����y!֔Hۥ����8_�t�]DB�MĜ����&�כ��ז{|U���
���^ ��$��8���S>��� �	��M�����.*m�[z��y�=�	|h�CG��Fd�Ue/�(�OU��5-��|v!��̸��q�v�_�D��K��!Oj�d;'�|�n��U�h�(I�S)��ހ#��P5
�2��)����n��[�V�շ�p���_H�x���j�nT�j��*���)�}�C&�����A������ҔߑJ�}%�����_a��c�T��G���%� x=�$�/F� �O�]�I(-J;�ҌS��~p����(P*�$]�2��l@Q�Jdo�3�G�����!��E'���W��� �f?��\����\p���>��fM�KF���JB{�8F�}ZW�8�����%$�9˃�(߆}o잚��=������U�`���( D�9���Wɀ@��309:���=`twB:�s��D�+ޗЬ5���5;�;ͩ���c�!�J��R����ww��q���ds�M�n�9�J��z���M�B��?�V����~M1?��'�E=� �cJx,�k�:�ˡ�}���O��ȃ�{)��.��(�Ip�[��n���i��rB�p���e�T��l]�x0��荧�����rܱ�y�ѯc#�� i}��7+^���XQ;bKܺh>�29����6�Ǌ�\eV)UPv�A����QY��V~��՗}�i���>���Q��!�5�D��3�5�p�P8���]�x{��i�[8��D�W�8���+�m�M)�O���I0�T�.�V��q�|՚p���@�ap !@�T���lp���� �![�`"�כ�u{����_��Py_أS2P�׃d�u��E�OQo4#��@#
�ap��NA{0�2 �mz=%��4���bU�Uu�n%pmQ��ܶ��� L�cHҒi��.$M��՛��[�V�9�����K��e̥�ZY����o��J�ĉP�P�a������^�k���<.Ո�M����0�^B�����T�+6�C]��,��E����g�*i�}�!Ȕ4*�޴��ɮ���Mr�38,��_ƞ87X�Sl�������q[�=�|'a�
p�5S����� u��hLGMH)�n@�)�h���#���X P!��~���-��;9M���kq�LR�Cg9�YFA!!�AQ7g��4�5_�Nj+�C8����s�
g�9���vQ�)��>���Ōc$G��v[2O�ʌ����j*^�n�;V���7=�D�U(v���K'��?y��;~X�2�fN|�ِ���N�d_�@�8ߡ��"v��>~�T*�ipvT�or%Ic)���º�O&�h<��|c�@RA�,�;�[�����ɩT�}&��>A\J?r���׬&�PC v����Z,l�Eֆ��t����Z*��G ,��fT�T2̒V����C�,Xܶ�rÑ-w;��	�Y��/xN�x�>!�ǟ1��h�I�k"Y�~<D ��igOv�Zo�^9�
�����S��Qf_ks���ؐ�C;yD���@zێvЂ��ī!�69��k��O�@�r��薓��)v�k+�Y���a�V��U�:/�@/�H,Ի�+�ؑЛ�FB�g`���-(Ĥ�C�pn|�{m(��aνl��B�p�o�V�}O~����*����ja���^\D=�j�<A�~��=�S���oSf�h^�Q���*E=x��Hap��ɚ��W��P��}�,�	�/�G�Z;W���K�o�j��z0
U˘r7���/ �6�s0�������!䖺����5��諏Ijw��� ��WT�2d��
�2��ϔ)��,�,�6h=�U�	{EK����S��g���N,���S�G�0�,Y���W�slV;�eR��I���*95����/\�d	x����D���/s��t^���-�=1�]��ѷU!]�������Z�iw��h

��YgmQؘc��1H��b�|E��b��q1,�[W���EX��@VBj�An�os��IV*�\��PہA9�ּ��`\ΧP�)���t����2���6�������pbx��Du2`�y��9sPSBy����͒3��@6gɱ����f뜌��(�ws�A���,�D� ��a����{qvx�
�^�t��	�%��]�!�l�82\6�
ʦ��}-�E�\䭖-�C�7J(����5\~�i�o.=�R�{ n�9���h��+q
�sP15H5�b	H��JϨ�A��
�Q4�&��}t���
t���^�T�V�=q0*�n�,� ��<�^�Fއ���1�DVw�o���t��H�e�I�)��)0��m4w����]��c���0&ܲ+e�(�N�"�"1��]FY�<�(�g�$�L�m��F��{A�	'���R�/��E,HH�x�D?�iզ"@bO��7ŀ2*I���ɚY=�]�����i��)*����w G9�*��WD�X� ϫ,Q�S#И3��ǭ�+�����gE.�j��;���W���^����ܼ��9�3�,w&,y�d��ʡ�d�I$�^f1�f �+	�:��O��1%�F�����"�V��O�1,�z1��|a�F/de>	�^��}��s�Iǽ�Ë�,���	g���'w˅3�C7�7PEyqz=�J]kx;�e]r$$v�%� �(g~j�e�ݫ�h���P7�bs��K�dF(�%�BItӮ�����=o��m�bD����:ð�r�=�Ym|��ٌ�7O��6�>���aq������2C��!yn
���H��g4�63u�r�®����p��&���b`p5}�:�K}�n�G�xսIs) ?�n�E�	hY��cT�S�E��{/=Е��&�},�!���&C����T�����u�`W�1����!���<�����O����t*P8��&��i��AKE�R��cRwɵ��r���Z���߭9v:n��T���/��	�eA�To0::��3F�ذ����������H�(��~Uɕ%ϧܰ1$d��'2}@T��`$͟���~���|~gU��d���E�W��y�����}kE���qb4n~Jg��8��ܤsl�R|�iH#��M��nJB�4�K��h��L���Q��K��� �#����Eh��L0��gEC��l-����5K��0��r���&P�Ֆ�	�F�Kp@[���;��r��'G���.����D��%�\?�j@���o��q�N
��eV��G���;0Y�������Q�޹�u�hWS�s\? �׼ja��	��]�u�~��H ����q��Z!�o2��_�l�X'+�c�{@m:{�@ó��_^�f5��e���edn���J*QQV'��r ��5+	>w�;@�d���Edf@l�?��BA�p�^����(��X��5��7�|�u M�|�wh#��n[��.�Ղ�ٍ;DG�����;���U(���W�|�6N֪�wk�(��bm��y������,Ғ��g�G���}�T���A`d�������A}���K���W���T�e戥Kx���ۄ�]�_x�YZϺ��DF�U^�Ӕ�،�-l�)��6�NN�U(i�Hc�Q�C�yݰ�0��A]�>���sj�Ȁv-'ė������;�p��y,X(M������n�����f�5>����P>h�]e--��p�3KG{}�͕��_Yg��f��Җ&��d[��T�h
�Da�e�@\(�M}9�"��q;���ò�[=Z���Aה���Y����i�!�0!��k�e�.T5lD��*�IQ�꜁G���P��N����hD�m���	pŒ#-~�)}�
+�E]BO�y�(ɼqb�9��9�z��u���������ó��t���欤de:�<��I�w���D�#��t���) �0��$�&
�T��-H��Z�f,t�Ԩ�:��&M>cU��JN�&�!��a�Vզn%����[)6�T8DZ&�"��ʗ�?��mS��y����P'��x��2.2�y���\�r�bWf#�{�\�.>���Oc�МF0���ڤ�'�Y'�!���\�_Y����aGٻ4^��A<J�������=�R��]�v���"� ���70!��l�Tifޓ&��.T�*��U�I������J�H���8������8��EԎ���b�����?fw�f�y�}!%K�]�.
�G���0 ��"�m&�ϫ�F"��Đ9l��̑��({�0�>��ubS���l�IJ�kޏn�!��؋HrR�YSF��C�8Wj>�lZM��������"�ڏ@�\�*YD����@�~�d-z)��-���E��~����Ow�9èG2���?n�C�.�ALN
*s��I7X���-�����Ah�I �a�*/�+|(T$�h��F_�+�'1�y:٤��Uz��l��*���ӆz-Ƹk"�
�n�`_%hSe��;��l&�U��խ*��B���k�Q"�\��Pa,�d��� 0��üKv(�/����87j�m�DfX��!��, ���nFկ�O�_̴5����/�\߻�
�P�\u���:������+ ��.Rw1��X��e����p���R̤��ة�`i#=�����Tq����_�5܂}a�_��fobFSE�ѝTvr�(%4�dY�Ԃ�*-2�p���k�%C�j&�T!�z�i��������ai[r �1T8����fC� Gd4�sтr7����0������T�f��G�$�~f%�X�(G]��m��|�U�v]�IC�!	�f��mK�^	�R��Ur��i��[2�|GG�u%t���O���wn��%�.����=��P� f)�F.*f�m���fz��觱��*��J�p��D�]�?����sa��]�ܣ�>��8&���	WB�����b%��9���������Bz��զ�w_�W��+j��Eyy�ۋn��Ú�e��?G�[Q��$���Ta�i:S%[��p8Hl-.�w�yT�/�9��g��i�|g*-t�*����i���M3"R�V{�nj%)�v&��ӓ�a\[;�2�)#5����̧y��L�+��& [��A�����g0�����|.��X��<*��&
�}j������=3$u��ʺ�������NAV���|b����7|���W�2�~�J�_��Jd��>�#��Vx��#�9�k#��Z�o��-�\�`��Ħڪp0����յu~j0�`e⼎�C�&4�ޜy��T�IYZ���dQb���o��Pҵԗ�H�)ͣI@=��"r�f�G���A(*uq���Y�u[�LzFD��u"n뻫6�QN�V��O�MFwS�[yk {)&��d������FX'G���z|�>𧺸�Ѫ8;�
�-B4Nsnx�A��� �sˤ�̵���`ֽ�U�	�|�V�!����m��w}����I�B#����Q�j��dʘ#���x���o�Sg���zJ���$��(�4�Q��)g��������b�a�A�A&ac:B�\k��2`VLp���c�� �F<*�Z ��(����3��>sG���'#N:�:��o��q� ���bOA=�iC�P��5���Y��u��ԏS��pP,w��ڥJ�Q�`yg��|]�7��c-z�'>\6�E(6�=4��F�X�� ֵ�H�Ի�'���Z�{>w&;\���Y�b�����[�ڀ)Ո[!��-h?�I���X|������[����x��6!�I�T �5����-y�N]�zX����\��Yz"A��L�0gl�ƚ�<v����d^4na2�^d��^�!�'�ҝ�[�ۥ���l\J`N����\�`mt���\�t�Kr��՝�y�z�2�j���;��Z��~s4�Еbi�)�/���Dvse�Tjc��y��5��"T%��K�M��k��'�,q���,�*eYq��z���yb_�(��~ʹ.�fʶ�Qy7]����#�1�+u٫Ė�lׯ%(�_.�;^H&�i�i(F����4��P(�n���mP����kφQ�^�서ǁ
�w����!g%�(EWf�|�z��2ϓ��H �hy��U=�\	l�K���	Շ򳀰���p�+�]BT�<��#F�w�?�������d$s0ի}c�#��بy�H�Q��R����;�{���OV���'�1��.�W"|�yÀ���o[6���Q��)�#K�R<��~�I���z$����`�	8m��3����\��p�JHjs��z�ޥ�W��}�`3�Č�v����u\z�F�\�s�t�F~U���'������E��>����fM	���'	d�l�p��/ORO�H!6�UAm"�^.�i�15N�X�<�i|�������<��~d@9-�\�
3^c��2�g; �k�}�g����7�C�~�\��V	�Sz}�����o�!�?�1m�j؃�k6S��%fį��������?Բ�YWf��N��v9{� ���Z�_^ 1!Ǔo��������k��*���.���_��{��+�5\�8��k]J���W�m-�^�4�y�nY��^�ȹ���PJB��6��>o��׵�V8pR�#��K"�m�X(<ڱ���X��@#�2���G_�q�D־!����/�FnA8��yR�^�rU� [�3��[u�;��06(kx�Y���R-{^�?`�
��*>�gf@�:&"�n�g��W�J1ip�6�ԂK$��I�[i���@�͹����3y�#�Y�;FPuD
d���⭽e.6+�8TU�m���0���à�����#���i<w0��]MGe�B!2�����)�pC�u�D�_����<�֋��\ɇŴ������9ų3�ʯ��4����ڌ'�۳��?���\�@Efa���98�$�czp��WNІ(���`����C�p�bo�A�豜D�c�Ujd��5]��K4�����@���*L\<�P\�0�za9;G��ေ4-���"Y��%��Z9���V�3�ΈS�-Z7П���H�=��i�2���Y��_�L�c�x�|�"6Bb[�Ov�iM���E��D=t|H�݂������U��D6Ʀ������"����s�/Q��Z�غc��3�SlS�匑`��R��Ue���/�=��Ћk�*DG�2�,#�sL.9'2�m�b5�#E/�!ט��g�y�π����GD?��¾�+�}��-Q�/&LS@�[}M�+?�nf��U��4�(�}n�r�!�H��j�'_~E�L�+�7z�@��˿_Υ�n��é���ؒ*�^ؚ9�/�8�~1��[F�ec�αID�va�t2!�S|B�z��-�Ț6ե����������f���Y�b��̉ד��L-����ޅ�U����v��1"��De���Z$�]k� D�`U+�B��\��흦�Y"]Ҵ+oCD(=���h���N�|O+�$���ų��v�P�Tc�`�=�+w8Ƥ��/���a�9������bD�T3�����f�+'dӽ�]1��8��Z���k]Ԉ�8���h7���bp���X5π��՞�pyK9����OS##�/��2��$g���\�@��*�.�ӊI9F���t��nM��ɵ���b��� ���	6��'�[�v.��6܇*� \��2�hu7�B��[�6�����9h�Ħ@i��ᦢV�jI�$��V��e@���)���*9/p_-��=lT\N���7g��5�����F0�y�%N3��[�a4{�JH�:��soU��M�9�w��k�e�D�3�b��F��Z ��7gc��8��Ӌ��+艡}�i{ap��-����:~5�N�D����n��y	�m��U�u.�JϢL��H����C���,J�s�b�wb=�AGϑ�E�c��R;����7ߓ 7U[?�Z	�iUq�ׂ���׽�dmWw�3i��_b�A
��}W*�y�2XJ�~D4���vWE}��p�i�!���w���8�m�W8���DΗ/���pT9��Y�P�?vWh�`l�@�_8�\/+�����\p5LQ�h��3mtěp[��oba��k��F��R�����~+�C�ӽ^������>�`rj�(w���d�8������I��i� �q���D�M��Za���C
�i���#;��Ex�{�9=c���Gn)�78�$��Tx��ؕM�R.�%!��]ӄe��xn�;�� �^wdR�\�Z���B���l�O	W��zL���ФY�= ����2eJ�g$T�z҆H1g8hJ�~ ޜ� ���l���*h�s�;�
����n`nش��}}q@#�Pt0�?��H����%R9�h�c� f�}s��o?���h.*Nml����ʼpt�1LVV�j�u2.�9��'ҫ����f.B�j�EI�+�u��F�y����5� �i��;��i 8���Z�g�%K��B�m�e��L��Q�E�Î���A�|-y+����Mv�:R{Gm�Ov�`^����P[��+R�q*S���2#��g�Q���WP�:`\k%�u@��Q~�ྋ4��{�7�bXQi�=�Y�''D�kǏ6L~�WH��m��T��	�*tkS �?(�I���.�6��Ғ��V�'5!��O(�s
�w�Efx~4)�Ճps��}Hy�vy����;#�9|�N�ըgG9�������i
5����,��TƋ?�D�o��TF+�5+�qS�ss8�X腏��~5�}>Ӡ�ӿ=����p�Ė~�˪d�κ������B�΢�4�����M)���q��m�R}7��á�w_� uN� �t�yJ�\(Z~T�͵��zs˜� ��N^I���hr���(7� �c`ĳQ�9���E�;��B������@�	�r�������}xv@�%jd����Tj�Xb��D嗫*I�@+��W�'�g�UW�T$0`uAR���������c7V"!A�9�A������/x�1���s�$-�[G-mh�#x����ZaDX}T�}E2x` 	����+���Zw{l�_�����|)���W�~M%�mePw�f)�2�mv�ɥ�^�d����xA��b��E�5q��9�@!�����g��U�We{m2��u"�0�S�@bU�lE����R��W���6���h�v�E5}����1%�&��jG3l opɬX��]X�s�Ѧ�gU �y]Whʽ�7ijs$��%��T|�}	4��7T������K~����Hq���8������ ��\мm����ä�:+�V�f���n��������1�N�^ ���H��ݤ#���f0�1?}��o� ��]f����?ז��iK�X�s X��
6������']��C~�L�
�-l�l՗��w>�iᴯwRlB���qp�1�GLI���CN��>�q��$����J��"Q�3\475�L�W�M9F����%vP��~���Ld��''�4���Y>�2����'>����A�A]ѭRi��x`��?K����8҄.���Έ��P�e���8�D�n��'�>2N���;�Օ�y�N����w�'�"����ES�2y�*��Y&��s��$7�FP�ԬMEG�� 5�Γ����ܦ�>s��Oj�Y���_�\�"F1\H�����c�ጹa����V_25xNm*
�U�L����vi�
v.Oacz���bt�����L�:��m����s�B�@�CP��n�="����;ϥ�y LM~�}`>7�=��(�?��G߰|ُ��#dE�),嫷`6�JFB�;!e@�?�NH���j���s �Ki���*�Z��~e���]q��#���������yS|c���!��)y�7"�C!��@s���&mA3{�i��L{�*��V�5���bap4�EW9P�-j�p�E{&]hһ8��h�NzG�ҏ�t��KN�E�bKY���Rߗ>�6�F.5έC�Y�4���� 7m-wR�ȴǣ=cp�g����FI�HB3E+�uu�AEQ��hDԘ�F���9*�Ms~2f���hM�uj�B�,�p��v�9j?$�|K;H�9����ECCPI^��wF���O�,U���7j����p'�Apt�v�{e�r�_Vw����:V��d�l��w��#�G�����K4�	�,y�%�o�37ZB���������X�gHIi[�����HÖ��Y���?�!���|n/S�ys� W3�k��SU5s�J�}��!�[�C	 �m�}Ģ/T�۵�\y�/g
�!��fĎ�h�-�"��.�1����6@�!���U�\��`"�j�ϸ__u�:6�KNa[{�/�������(�=LW]�N^H��|�8Ա�U�)�&�Xy��+����_��)$��#�'� B%�8}w��.���d��&��}��~u�Nu^�\�!���m���H7}�QT�#�ܨ3`�0�qy�^.g+�^�+�L�a���ę�XmS�z_@UP�e���j�6�/t��>��R�o7+��ٯ��3<�2��b���hy�=��4ѩdW=s�I�j\�r�'�E�D���m�#�,�z`�ױ�3_E:���}e��/GBח���]�K���mDN��55۝���S�
A�^t%?���6B6W��n��ɴ�^.ɾMFW��-�L׿C�ց��OC��g�� Q�N�Q��4�MOW��d���\[�q�{�;��LԢŤ�DW��	#q��Ɲ[�d����ȧ�~�)�2�r-σ�"��~C�����6}ԽA�`?�;���r�f�@����/�L9-�?+v�oX�VR� AXS䣞	�z����g&Nv�[sw9�Ǣ��х����QvQ����9ޓ7�IV}n���Cg舻Sy۞����6�qkչ��7�!��Cӆ���j�M5���SmѥcZ<1d�mW��$?�aV���D΍d!|:??@ҍ(T�-B��+��aDK�!�=�<�{v]8����jo�Y�����Qs��%�Q�kw~������Jd������*P[�0�w��c��`vΗ����4)C���&,>����`�;�0q���6�$5��EK�dNS�jM��X�Dj��,�L&�Չۍ&�E�O������+r�3T�$�$��^�I���4�܃y/�>�	��s���!��b�AL�uh�2R���yvQpRx	P�}�إ��CD��+]v���_�U]���7x�f֫��D=�W�E�|ۄ�,�p��[v�]�d�d�\��W�P�C�%~�A�G���LP �4����UG�/�����ހ��1"*��9�~-?�\�v �|���`��T��ɍ��?�d����wCyhf��*>��M�s�%p������g��;A�{z葔ă�U�d(%�Ө圵�rS:�~*dZ0\�}>,��������[�)��T�(TY�M���P"ϪE�O���ԍ�WVE(�+�X�����}��F�p��Xk ���r�h��Q���+D���:\\�cMk'M�s&��lڹc��#c\^8VAv�P#^R�����$��q���%����Z����3���7�l���.����TM6�)W���4z14��[X�`O^�������SJ��^_�X��r�V�~�=���s3Ǟ�6�E3a�jd�j�M��D��#�`�.��ֱ+;���d�
�jqfh߉b��v��E��F�Q�����M�=��Ƌ��<��E��>goƴ�Z�V*ߌ���e��qH������wf�,es��W�����E����e��v��c7�����;���w���n�Ӽ�w�Or~���Ĝ����}���Gi|e
W��@�y��.Ђ7�N�-��}��u��[2���{�
��Y�@�
BF�Q��d����<a��������?Mr(����F�3h�x<�d5�硫��tw]�y9[�G�sfY"��9�B<tTi����Na<B�?}4�]�RH�+�7���]��8Lae������Iw%�/��x6���af�u(�`�k]������C�}b���A)#�{�gĢ�|��p_���VjNUO-����'!�ǈ��|N��!���LO�	�ʪ<:����&@��:8�R|inmL�q��uXv�ĸ�M|�F�{�Ǜq<�-YU�#�BB�������sE��c�����x�?ׅ�q���$��p ���čf���k�LCE��u�X�
��DfSp�/�HSC`wKQʌ7b���I'%��؉k	��S/W���p[r��������i<�HVI������qn���9�f[�P��N�>+���'H��d��fOZ�җ�~ ���n̓x)'�m��G	L77>�����H��c�q��v�0l!��7��4�ե���J��j)$��7GvWm�Q�|���lS����-Jv�WƂT@�(�qY�,�B(�ߵ��ErʘF�ݳ/���,Y	Sx2W���2��#S�7��!�(ԯ��3U�Q��A0>�櫈��#/�!���ࢉ�U����'��M��q�B�����'�yB�IeH���I`Y�-��r{^�w�[�!0�Ӽ	Ʒ�ق�FA��eƸ��j���n���(DN��=�J��a�7������M��w�Ҁ�M8z
7�z0���S��$|��u�e��za�#Ԩ��H:�	��{����y��̏��{�w���
H��T����ɮ����İ��2��W�@�͊������<ǈ�B4v�z��?�Q[��z~ϫ��6��� �ߴ�UC��n��khs2;�X"	Ơ0�.���(2ˢJ�iz���T�ǎ.�\�BRb��)������s��ZyH��o�2e��<\ςT��*�.�SU�����#��H¯���b�_PU�g�J��q�c���p6 �_.�HTwsF	�K���(�<�-"26���� ��q<���C�̞����4K����JҜ��R�i֥��=T!0�u�3e	�edx�d�O�����0b�#���*O��i���حvZ m��y�l�Ȏ�GF�*O����O����)ո���وy�&pC���.)h)��ީ��v���_�q�s1E����bW��m7�!DP����*�M�[m������`�,G8���B���S�f/�u����:V?j�l^%��uM:�۔��Ò�0	�Bd��s�n ۳�w�Ѣ��d�nfIƨ���x{暮z6������=�8�{���f9��X4%�4[��z�w������}(5��)铃n�I3(��m��{�jП��ЬF� �׶�x�E���)�"���`���D��]M�6�����l�"
S�V����Ul+��\���s�1�5Y.���0+���|p�)���:��6+�t��:ėPq3&W;��P�ݹ���6ү�*\�o݈�u��xY׭)밻i�C�!y�t"��ܓ2��4js_*A���>�%{؂%*N>��#�jw��*�Ζ���W�^��E�+@�����x��� ��H�Ֆ$J�21��:���<�0�����t,�#���J�i��� DK�g��*�/�,��!6�)�#��.��5�O��"//3�2��@�t�x×7�BJ;r۷y��
��!�h*�*�i��o�oaa�o��O��1��|+.Ԣ���Y?&7.;��[L�r�Ԓ^
��1��W[R��\���a��k�F��ٙ|D����f+��jM��2ɼ��L���~���ZA[��B?��h���fs �c�]^7,�^�D�.�TûyŒw㦢�JL=��d;�c���!�?��W��ƑNn�ʢ����)F E8# .��3��u:��ڲn������b'�SO3�8P\�Gg��ʤD�����E�gu0��QI�VL�ѧ�ǘ�ax���:B�W���;��=�p�g?�>��m��j5���"R���\�7�F/*����XI�o⓱�d9���.2b��~�,�D�(���\*"<���I����s��g�U\�$�����ϩ>Gr�zb?A#��t&��ia"0C�y-��ؓ���'҉r
8���Z�hc�4;�QX����M�jW���o�p�Y�㚝f�[7z<��Wm�R�����}��T�6�#�zk��vLӺS�M��<~F����H���X�?��d��3EN�J��衞~lOb�[�u6��H{����I�
�B��x���u��9�IKM�y\ ����Ǻ�+�ҎU�/�0�� ������|�>��-z䲃��б�Ԉ��.�N3�@��W񺙫���3� �bJD�, �j�;9�*9��l=�īm�L��ן���~C�C{��a�3��H�-;�[@2���٭ �a\��R3�4����qUw�lA�����V0Te�`��?�l�� �*�Ƌc���ﬞ	d�%���bn��ş�Ⱦ
���;Uf>o����A��W��}��G��J�BK��b���mX`��<g8.�c;��7Jc��
�.	۳��Kґ�Ь�A�+��V�&�'�d��d1�f�g�ɰ�e��� m����ڢ�ꑯd��BxO�������\�΀_{Y�I�)(��w�F j��W�z�*ϝ�G5�l
d��&���;�8�3�A5�Gy�nKT�e`g��h����j�)U�2�g�삸��Pt�A��z��p��xfx�%��ߴ�	���Kư&�yyO "�������n;F(潹�D�lh��I8�~��������՛bVq��z�2حǝp�f_��F��>-֗F�n�L�3D ���<4 {4���O���+҈�U�8 �����A�Y��T��Ǯ��'	�c��+�M�1��3�rK�(����Ʉ���'���CQI�*}7}74q����6~E��P��o/q�oa.��A5㙛I��Հ���ɪ�z�ۂi^ �=�v���y�����S�A�t��Ϝ���).̭r^�|��;�hKBM\�j��4&���~!l9��!�4�$�ͷT��
�J�����u9@7�ue�I-PH��gV�,8+���������F��@���H*1U�}�"i��g-C����&�!��[mm#�t��+[(�p���?SLB���2���;�b�n�El�A�[��"|�Qz�b�SQr��e�Aj|�d�����܅K�z���lo�s�T�v���������~|��x���nd ��P�@2����������d�F��b^*�*�B2`�F��/�zM.�r�Q�)~���t�K<ɾʗz�=3�mm�ي�� b�I��$�K�
G��"_]�_8; /fZ�η:"z�)�Kg;H	1�6F
�{n����(̎P}������5��L;��57��HM� SW4�<%l��
�V(N[<��n�9��7���1���6�oW�L�1���W�*�x�e~�hs��\��t�_�f3�J�"&|�{G�C ��OI����	Q�>�Ļ�Hg�"��KX 
�L��bm��½KS]|��N�G��C����H�?6uJ6�lh��Ho#)c��()�iM�_=*�\)Dډ9��9��j��Q�4��d_�q�t� %�k�_)������{$��0�p[؜DD]�ڟ9)N݁�r@F}�N�"�k�x�_��ZpQ�oϠ�O�s{D���t�|o4@�Mc��쭨�Ǿ��Mt���E��daX�Z���G�$� �j(�o\�Qj[�Qg������؍��a;ǌ+�g/�� �����Es������P����hV3�9"��i���p=�j,����1sna��v�$Y��A	�'C^J�4�&o#�oÑi������2��*}�X4iU��Ko��p��w�����ps�؁�'��_�����(���>��{��&m0t�#샓;HړIQa��n�{sڴ���䃌I��(���a|̀�"�2)h�Ƹ�#�|�B_�����w��J��UWqT���_��v��+�����W@�z[rJ���O����%@�Gi��言��t��]�Yv&T����q����9@-zy4h�VۛrccNb{�;���L�\MBҿs/!HE��J��+�2�t�ڿ�B�p��]pXJ�*V
RW-0��ښ�^�إ��WY�s���:-���b�kA��
��n�j�S<*�(O&o��Z��)�3E=X����1*mPU���uS�vvid���L�2�@����yQ$4�=ݞ��bIwQS	>K�?�9l�����*8�z�1��,n���²�n~=�dٷ�&}i�pv�0q�8����T�l	M	��l4��b�r��n=�R�\��X�f���$��xW5!�3fr:�U�'v�C���J��Zo[,��<T*��WE���t$��/�u&�e}����R�m�¬�3��Wu�+�9n:\��v�	����^� �$�����t0�C�A1�V|g�.os֌�{;p((�:���La:b�>,���y�yy��%�J0/��v�!ִj<�F��6���Q{1"�����Uc'%��+�=��"/��4�<I��`<=��ˈK`f��t_����T�y�c�8ZO,��Z|��1u/��
�.liV��8���Y��� >z��<+��X ���W�q���{�rcc��l��n���m��[���r����"߻+y ��N��ȴ '�_Z������U������jl �hP�˭A,���s�2A�oGM2O[4�>v/��GZ;���7 �}h��������Ћ�[y_��bwN9�ֲ��u%w\�n񰄡ٹ��R��lD��y[!���ky�Zӝ�}��Ŀ�l�F�V��!VdVI��ÿC�����]lѬ�E��o�����E�e�+�Ru��������`c���QHج�`5K�D}u�у����!���N��^���N]"�Y�4:I<�L�(�u{��g�P�Cߴ�fF|��Y�g��*'��F\�W#;W4�JſpR��Cۆ!�����(�a�9��_�0����>a-=��K��)����L$���6�~���^�%����1��)��[�?_�8��Zb��@��..IZ���rr���/����۠ �W�y7DǌD�ك��9�͵��aq^7E�xf�BQ�L��K�> �+!������x���~�t�|_�t�14�sH!��羧$����t[]M�;�y���`6y+ieX�=.�2���Oß(�DyP��+F�ݽ"�70���t�5�@�DG,NQW��D��Y]*nQ
�ې�@��ԧ�\�����_ѣr��b�gEJǠ�u���e	X�wS1�Blq�z}�m���#V�=� �-%ܳϔ�;���l]��E}�Q�E�^����_%Y���2�
�S �}yb�P~d�Q! \^�d���ܯ>[ނ��<��/������d����EA�m��6>ê�e�!e�F����Q�$��ա������2�����{�$h�EtX��TWӹf�E�e��kިr��_�������M̩8�]����V4��m���)�����_�.�w�@t�+�S�j#' m��`}���H��u�C��.��#Np	?�"&R�H�p��YB��v_�y�����8�1N&�d�E� Y�F�琉1 �:1r	n`��������@\�L�ߐ)%�����3����b��|Li;�%��ݔvH`,تj�(��S�}�f��*��S(��]3`W��k�hm�����%/wQĜ�!��bs���~�¿T�,��n�[����>�2��x��i�Fn�e��c��֤��\�NO?&�{�{����aq���w����Wu�R�ۗ�����CԚ�R�QU�Ic����~	�n�>`���5����ڏ��$վ#�����H֖�|H��=v��{68����T���h$B
[�Ȝ�k�υJ6��_�� U5���JDR��]̾��$�`o`�ji3�E^鉵�N����?C����_�	�Gw��w]@p�ch}���5��:EuB�i�� ��U����,��K�E���'�4�9UAK���*y"�!R��+6�ə��}N��/i\�����%�wYe�z����r�NX�ލ@��_=��O���A�Lf0�^��PAj��hպϬd��*���*��Y�az����"_��;D�H7����{MV	�S�@�΄}���H*y�Ո����/��m�E��m��4Y�	�A������u��,�:�.�:��D��+5z ������j!��� ���Io^{��ê�Y)B�,���o{<���8��/�����u�ܝ���N
������+�|C ɒ{23�N*�RDUL�5Y�	U,:�:���]�������9� 9�\s�C4׎B�+�q������z:����4�>�~�Ν������[�E��7@�qʡ�ð���m�]���|�������5�(cY-Q�>�Si}݇C+���.aw����+R�ù|n�w���n �2i���B�mt�����٣x;��C�߮��QV^bFP�ʛ�.��jo�d�1�<}zn� A�F:9��G*i�J�� �7�4�O������d 4��k� vqH��Iu�b�+'�W*�!�ĉw�W�קT���*�OO�+7x���,�|�*�r9E��=�,Lu�2���j;�d�ׄ:�zh��{�d'ܵ{"���8�a�2J���jG��D���m7ɺw�S�.0A{�����!��Tl�OS-UlD���y���j�Z�i]�w����b�$�9�����!����C�:�б c���peF��>V5Ť:t�<&lJ��ǐ�)�6�̈��9�{I�k��l\~�gnX�܊j�KJ����8E��<���k�H���S�b-Z^D�u�_���I'��v���q�h�~�R�ys� Ƶʺ]�c���*N�6��C#��I��f�k�r�d�nW%�ř��(�s�N���=:�G`�Z�Ń��fMw�c�:�va����R텖~�\��T�EH~�Q�0�<���z�ߋ��^��ڊ:����\��j� �s��)�/i��"5ܫ��9O��Ф%l��J�s(�6���$�}=�_�m��K7t;K~[���g��S���� `��┿G*g]~d�5m�fyi�����G�rj
t�4�	�	)AS�T:Ýt�A"�/h>n��D�9~�������|fP���i��]�W�h�Me�����I�]Ձ�t�B��by�q9"+x\��h���w��+5� �ze�E^uD�����ut�68�R��J���E6���`��w ""�	hYQen��DuQ9���uZ7+�����AFw�X7����2n������d.d���p|���#���&���;���"E[����j)1����NBUo\��V��Lt6Cei��MpHQ.���vtaD�^S#��tE���Y�$nF��t�UT�ğF�^v��b6ȇ�F�5��J���	v�/���Š?Aͬ���K*xjfm�oo�vՋ��cGWb{b�`�f�h�u�z7>Ąc�q�0�a�Ŧ������9C`�P���t>���b��.U�d���wBXL���m�ov��ƱJ�V�V�r���}D�/@�5������%0�]VޓN��_����R��F�r�y�r���ݢ���[�jp�0����LwC��*��95̘^}����E�f���n��O<
L��e>�ab�K�by7VF*W���$�@��7C=!Z���K�f�6+����m�!H�q$�&�TJ�I�d��q��rﮈ��	L��͖������J��X0���6uZ�?��]�z8�m:�����A���d�Z2�kX:� �B!�����/Mr,1�O�>T� s]h���Ϡ����E�&�?��d0��^�ktz!���opΏ�?0��Lq�f��ᒠ����ݪ�J��w͎��_���[���eP���/VZn�>ϫ|��t��EH��D��-l%�#�y��ۨ��96v����Z=�Ȋ!�<�`T�ˋ�+�(��g"��)�`N�.g�W+�9}�(��g�v���]��2s�q�L�s�x�*���8��msvUiX��q8����i�G4�����;���x�	���)A���yTNf�La�&���^�0z��g��W���u�2A.P�P��	,PAE�i��k�:}����y�4Eh�PX��<��`�������7�[P�I�����|�Q�l6B%��'�*�暕�8�O��K�&�����^�������>���5^���av�v��躪��A�W�|R3�
%����j���������)z��1�;�A+[=I�:���DR|�3���}pAm	"ޟ�f&7d�����&J)�u?T)n�U�G�(~��;����C�p@�N~.��=N�jd�3Lk��L=]n� [-3���Y�1M��zs|?8��х��ec�Ă	P�P�-	/�vb �l�&S
g�7O�4�C�D�zWLִ������%�G�l�*s���ɋz6��&��K(ݵ��[�^��<�e��PY�W�C$n죍���
���]�|��T	wR�]RNν�I��b҅�ѱ�x��b��$������x��<����\�� 5�S��;Qpv�i8�c����6�����oG��k��s��Ef�E�=C��KN{�m�f�:�J�]�}�:��$�TIԹ&<��!'G�\w�J�H��O��J�9\��z�!����}�ٵIs8�4��*K"�hL��e�F���U%�@��C����`b� ��˫X��v�Q�x�HI�__X��>�<�^r!���EN&��E\M��C.I�	� ��v�)K]����p���I�5r�3�T|�7�{�|a�I��sC݃?`_��_ڎÞA��73��1HZ\%-��(��a^9�n߃���-��\�0���%�3�`i�y���Y��xU�<��w���A��}@��U��,�}�x�²R���s��͓�ݣt����qvmކ��Ԝ�=��߃����$C�ݜء�� F��8 !�������\�1�Œ ��#���Q���R���/�qV�w���HV�7�9L�BՏ��vzS��y������<ʱ���HC�x�Jl~���8��"Un<]j�6LD���Ƶo�������-��8�����ӟL�b:F�/�I�o���,x����q��r�j�15��$�SI	�^ oe��!�y��Э���`򦚏d�,l��9]֮a)�3�&��W�?�����VO+��Χ�~<���f�!�I�M�?7��p�ON�+���>��oENE�v����'1�d����Ғ N�g�.m�)"��,� ���vޒD���=(R��r�&GD7�>O�!��e�l3���D���~<ʏl>_�C<5�fJM�g�rZ9m
����f�0�r)�@���B���Y��x��YȄrt�;k�k9�����4L+�ۋ�P�]N?C��)���q&@��F���I���;��q*�)��4����N��iCp&-^u[_
���o]�'��P�(2]�B�"��i �s�*�����&�f�@6��
)�~�8�<L#o���שE�7�F�udA�����61�r��rֽ߶dHv_ۜ�@/�8�E�@G�%3J�z!�n����+��}~o����)�ޙ���9k��������܁(�ۗ[�,�>����R,;x:��&����~s�@���(�`�Q��5� .-7����ĝ��5+�p1�}$N,S�"F��19_��	*���k�?�������;7���{d5h�d6,����hut�ef�����X��Ht���z���$���`�'h�e���ā�Z]��A�C���AJ4Ʃ]�M�����`��٢+�_���C@?���)���o
�pp�ߔ@y,�*ޱ�UU�Y3�[4�<�&k���T�؃���B�y�fW�vA�wJ���q�`�w�Lms;��t�2(�G�7���O>�>b���4+'�Gl1���Ș��m��##$�L�п�!�*�y��~�Il�x�o����)�T�J	�L3�[`p~��6HT���X���ݚ�z�\�\���1J<3h�9��&UXp�"
�g̟��{)K�l�L4m�lC��q�E�I����cB(���hZ��-�J+H���X�0s�-���<#�~6��xnG>L�t���4Zk;��A�}nh���l)e���_lae�y�7�$H���q1
�L��n��>r��D�����Q�E�ԭ���1��.n>�ҕ�b��Й�^/#
gUL_5k@�dЀ�}��Cϳ���O�k�� ;\Ʒ^-탒}�F:S'��iy�>�b�_�#3ŭ���=8�jFڛ�濑���,j����+��&���φ��9{4d�Lk!.M(6Lkx��uՍ���*�iμ��R�P�p7p3�:���.Y8� 1k��x\�g�'��("|��^�T��y#~3�6��3m6ϊ9l���)v��>f�5�y��Ł����T6��F����;���Th�i����
�>���M,M�S�E�-�|*�#/ݿ%�������������LS 9�Q~U�ǘ��s#D���x�S���������}�)�p:�B������{^@
<?݀��{h�T� Y~浥�:�>��]�߁E�aA 't/dJ:{�?I�A~`iV�pY����{�_|�uz�*�O�����y_N��z���uT���4�R����C�@�r�w���n���@a�v'r�*��?����m���r��f.�;�̎�Q`~X�l@��"��A�j�R��$9t
I��_��j�޺���������_s�}�cȯ�R����;L>�G�y�<�7ؽ�z�#Z���ʝ��ߙQb�t�Ʃ��y�Sd�$f.�I�B[0�-�2O���T����] .������	�)[.���Yk��R���.����Dx]�vf�������_A쟬���eX�R���IF	g�������6�T�?�8���F�v��Eh����������߫0J�݊7OU�G�|����7M�����|'HzJZB�&1B���+m��ci���;J���PE.���]M��;xU5���}�l���^�~��č(����]I��x�z�aJ^0��������޿�l�����s4�����&��ֈy.V��x������H�2�۝������Lig���b�Y3>qY�p�sm-�n�r1�\�￴�� �{���Dl��.���;4F��ġʯ��hߒ2o�{�(D�O���RV���k��Mѭ� )��j�N V������C�7$#�E1��~|qI"��5&�`�Đk����NN:�nX����������Y�_�;`�/*������X�!�M�ع� uB{
w���p��I�r��������ċBg�����l�ͼ�&���Q
�h��>�gHr-���8�N��a���j��H��W����W3���A�	ǐg �۫���p(E�L����|��ˁٗ��y����W(��?*�����C�v��ި�@#=��FS�6q6���(�.�z��=���g	~�l�4C�6Fs ���;ڦ��{|�i���v�i{	�]d[X�����g�9�ߤ>9�iW�vk��v��ǝ,7��U�(��Z84�d�w�cB#g���:ZߵƝ'�?���D��)�A¾	�rʙ�*���{��+.ɢ8�7�G~EYQ+'�H�e+��h{ϴ��E�H%��Ό7� kZ�G����#p���+v?$�l,$P��₹�()D��������)��#��Xa�Ư{I�wmbTU�0!���D,_/��,��
)��Ħ��:$�u=H����~���s����
��I�Ȝ3���yD���F��^�w�}o�b�8VK{u�V�(�?6;ƩZ� ���Z��	��(U��ތ2��W/ǬNy|c/}���JӴF%�,�l �?xr�6^���e마�İtskFe�il�)���߶8� .)Np�"$��A���G�yLr�5�:E�=��l#0rf��7ކEE�t�X�8����GP-��$_��nTp��o�<����Q��D�W���lM;���{])c��e[��V���Qy7��<�8����{�f�3BUNwN$���.��~����%H��n�N0��' �B�3� x��G����mB,�k�7��m��B<��b��}|h�>��Ji	����Je�OS�xi����K�2�[m�K��-�ˡ�����k �8��I���oF���n�b�g�[�b=��(�+Lg�.��X�A�ʎ�ڌ4���#No�N�]��;%����*�]#�caI�������E�f�vh�t9���E����⣔ 8$�
h�s75�2~C����D[��x����aV�|�{�.���%�&([B�&s�B̒�٩�h�o�m��
rp�M��|j�C��q|�p�j��:9�Wr�~��6���fNQ�z���䎭c$�oر>���i��cw�:��
UB�8;���?S�Q�q����G?B�iض����z���T¥a�u��s��쫣wĮUG}-��e����h�Z�"��d�6�@"+o��B�5r��t��1ٕ(W�}�Boa��U�y��Zx�F���s^����A�^_�` ���X|��5tB�+��y�� ���=� Tz13�D,6X`�g���a���K�[OS������IRf�O�V�K�cn���%���VJ�0ɢ��P!
�u��<�s�������,���v�r-�?L���]3�m�lS$����4Q�EVo���oY��07'|,�����V��@X�$)A4;]RR�r5��o;�"�}�uءi�f��^�_��~�9U��W���B��n����K��֢����{���e�b��-`C�p��m�a���&��Ԯ����|�#��T�(��CJ�$����6N:��b�Q�n\�������_�E��l�[�N`"k߬3WQl�tM礡��L�wV���*۪��fΎZDć���� �5�#�އG�NQ4KQ2����e��͎wC>�"9�����Z�ߢ��y,�jF)��f8��Z�TZ�GCi�u�^Ѥp�Ct�E��m���?Efߒ[d�QvI�#��9�����5>L���jgW�r��D��!h�\\���)m!�R�h��D��` ���{��a���E�w��r�$H�4b����۸�煻�Bn�Y��A�g:���Vɩy�Y��U��3��;g��i�!�1���ݭ��X,�eS"ߎ`�k ,��tԋ��N�H+"���s�x<!9θ��{ �%G�xY�%�O.�<a�Mc���գ��[h�Q�gr�k���<��C���y�\!�#l\�:�F�˖�&�M�ԃ"���r@˪w1�Q"Q/�`�3GJ� ��f�e����R,�W.��%��lۯ��pu��@u����hPU�;�Fp�uy��?}���vg�Ꮆ������:��L/|��B�ٔ�)rSs�����\��������N^�-�m.z�;�����֫��|��y��j����8g���ּ��qXw�8Ǭ����s��4�h�&.t?��es�[(��Լ���F��P�>��f������޵@
MTg�7�&�ѳ������f6ϼ[y�͍�3�F��${U�0��B!:��+W�"�jg��h+RSL�����Gҭ�x.�^���H��{�o��=��'2�xG-z�G�v����q��g2�o8�<�E�2>CR�ɶ��U�IF���Z�Lɕ�-UY�!iQ =�@n��Bs� /�Z�Ɩ��xlY�����x�]����(1�P�ߠ�<I�W��j2P���OGF��$C#��b)��84ب�e��eA��&�1�2g||c�`ы��`�\�f��Wh��
S�e� �`�4��`��;�!�3+�Q=��9Cv�@� �k�DNLɗ\�m�.���T�[�_S�B6EЖ[���M�n���fa��Y<�&6$�ؒ���1ɗU'�doU�J���؋@�!�z�l�,oL7�J�"���j���̠�OТ��V	d�h�,O7���	#����U��9nT<k"@�dC]��=��vs����8���]3�73����r��@0���{ø��Fb�Q���	
�c �52��+s���v�}��o:��*1y~t%s�a�Z��<gc�ު��wYi$f�ǐ/ѳJR�̩�����8~���G>�JuO&���5��Q�Eb����zSaq��X:1r6��Bi:A �����u��N�*�*���ı�g�ɲ���b��{W��7�,=D��	��r��К�l����^�&q���śf������y	���BM�ܳАMp��-��6ވy�s3�.���4�R�+܏�c�&�4��ig����^P��B��I?a2��
�	AI$B�#�����T��\�U~�<�軨�Y2|!�ڻ)����z�������ƿ2h�!ո69H��k�da&2qRzؓ�����,��շƺ�bM2��L�߹Ĩ���\��o=v����a��q�8�gj�'�v�v���˶�i�V5Z���!�<�c�����n'�x�K$^��'�[��ïi�uto�a�,�UEr��P35��s3���p�
h���9����/���>Kd��Rir����M��Y�������v������J�a�ʈ��`T�vr�� �Z�$p�8������e)@�Y!!"1����O��ue��>�t�t0B
꺫�m	���cH��x��S����bt%������eY�/�$�������D8[m�foD.A�9���R�˲!��|��>�Z5���f������3��ļ�B����3Q���τL�Hȗ�C��e����DCw������<4�]�&Y�[�R@�n/.k�a��jthU�����J	�Q^#���_<�W�ڰ�_@�
A� ��!����D:��h��C��~cHӧcK��.���V�d'�'�&��zF�#�J#u�n��P�r��jD��4�w�e��)f��U/0��ʛʽh6�8Mq�Ρ%�7$��h�Id[�E��f� ��2��g�4�0�}�X��ʈ�ǣ7[�_�QA�]�派m�1��<cS���?�.֌!�������Wm�؟��?]U���붿%n������ܠSz^�}w�}Nz��10�-f�=�D:�Xo�P7o��!��ß5�qn��>�
�]�#����DUh�ccvm��d�T� ��:����.�vZא�y/�0s$H���5��4j/�hYn�Z��'!UV�7�~���3b�� ��䠸۔������^��z���c,�� ��m��.�d#�SX�KUs��eV�+���9b-���g쒰}�]�_}�Ϫ�ֶ��V1�6��z�	��g+(�����|�r��c��e7���{����+C>{ ��w�@E_�wHa�RAn�Ĥ�y6���6����Y����,��v]�0N������V���-�mV�c��9�eމR;�r75mh�"h���Vig2��D�8@�ײ|R��m@�z��KBz�fb;h�+��K�g��L�?��/L�1}?��`�*T}�&�xT�;��?���4vIד�$h����r�7輿<Y�^v�B����A	y�6�W�9���ߌQ"����4����Ek\����i
���p�E����j:v�U*�Yt�����a�ڱ#\Ys�Q��xNv��N,�d��G��a�̐��n^��w�����ֻ\�5���뗄[��L�+>ȁKZBRn��)�9���B�H)�� )=����}�!�U��*N���������^D����Q��r�v+�+L�O�$���\�k+����C��>˦dǞ*C��ᯧD�!�xs	{A8�+9�6?�3�J>�c��G���8|�@�j���c�\�1a�� ���s��ձ�%���NM���v0�"�ĥ�rRG��n��w�'1"�\E�v�����e ���Q��z͆�W[�� !���� 8;7@�j.����� �3k��>�����V#�CG�д�i�I�A����<0C|@,oZ3���wū1����{��5��j:��i?A�l��8��=�cB���6��w�A�?� �Ov��� �c���ye���w�.���<��M�7��-����]竟D�}�GW6闲�q����F?��\my�(�\�W�ٟF�Zx-�ibXe)bs��|����� ����a�N����_�~Dy��}�!<?X��r�¥v`1�a[�S��C���|��M�-&�r/?Y������?.�E��tg�?��B�_Z'�.�g��GF�d7��RHh��&<��;�[��_�?85g�BV�S،|�c/
h�9^m=OQ�����g�$*���I�r�#G�W�]�!<z�`��"ue{�O±��7���!��?�	���w��!a��;���^}��U��������B����ޓ(8�9պ bY���RS�%���x����ig��U;� ���f�	h�� �v^�"�@���B�d1����{�G}�k�S��Wb�@ٸ0�DGЪ�={1����<@D
�A9b&�
"�eJ�~&�'��@F�'#Hr�tW](�>�����o���uf>���z �����,"�E�(]571���8�X��#�!��i��2t��M{��ꄲ�٠�P�[�N#��f�N�\ 9_��6��,l� �,`+LVWd�I��q�79oo5���bC!u�9k�ٕ�]љ�]�PBwk����1j����i��M�����w�;�,�X����Y�t��+�V=��A	'��M%�~�T
�f���d���2�!�"��ЖY��J��S�f��
�]�����\mX��7d�Ȓ�PCJ͙/��5�����}[�z�(��G�d9S��4~���fT��1y�IQ�S�>8� }]pҌ|w(2��~�@���j��~м�`pfuh��~�(}��a4\���u`�H�w`��ڍ��˞�ed��{�?����i���?��1B�ݵ�I�� ���m8��uʮ�t��U|��tL�J���c�l��9�
��� n�Sleҝ���T���qJ%�D͌�{`������K���|�FZ��_���r9��.�>�gy8����mx��	�T8�U���-#!干�5���䊚!���?�@ e�ixώS��|TѲ�J$I
����" ]�!@���n�@~P��[�0��w�����Vmh�ͱ1�<sk;4?�����_m���0nY��
�/hnyc��?\�4J̮9��W��f�6P(�df,"�?�0���YX3-�q����>�"����!�ݹܤ!R�]	g�D[�nD�J�#0�bL����zkx�	�D�`���:�hZ�v+�|#ni<8�nw�� p��e����]�H"����͢�/�Om�f�0�EXǠ������kx3mԜ�)rw�$�1ӱ�2��(a����]ǲDY�2�w�B4���@��w���',���-�� �"��b._X߬���hi���:���Q�������C�߈��WH����ц�����@L����)2�F��t�z}t��]����s��y��'�rMC5�Ş����OK./L�g����u��Ȓ[��tRqO�ݶ
��x�<�R^��v���|@�]�B�����Ј����������ל����#�ms+G?w�Z�j5�uЕn��2����/�2�y'�~Q��7��uO����J�q"˦&�YmM�#���M�h��K
�VER���{���V������R�@t-y����<hۻ���Z����ۭj��j{���RD���ј�J�3#��8����wU�lN�N�	%����Ub�M6ʀ7�ZC[^�xx�hD��T}H����9�b$��)J��r�6�</h� ���,ĸ����'F��-?ӥ~��S���U��þ��/t��2�u.�T$S��CD������R_�?_P��k�I�����L����� ��<<#���So_g�]3�ަ��U\lT��t%bN)Ν=f{�B�Lk�h��c��ֳ��S��a��C:�ُ�Z���6n"&� ^�1���]��VЉ_JP��z�Hb���Sی�y��h�ܛ,"�E�L�$)�0<�Ԓ֎0��� ���ӽ�x.�定9@�s�uϚ&V��+�����g�|"�Պc� 9�z�xAHĜI�rٲIJ^v�g\ �{��D�+���4�*:&�2-��;�%��U��k�$�ڨ#�3��h���Yt�V�T�Y9��r��b�|��se�(=%��y�:A[-v$�� k�1Pͺ�2X%�1?��XY:�ݱ�?�p)���%_!�9.F�$���H/?����d{�\?h�.�'�Ͷ�eGAYU��df�-�ؤ{rOZI"��,=��r�-vXl��E��ae�r��E�հ��С��G����G�@��&ת���_xA\dpR����2� ��3�����afb)�4j6��E���`��Z��9׏�(���"�'���;i��O~���f�i�y}�������@�ͺ~0oTS�3�#Q��<�Q���v�x��@{o�2)�<)�b����A�1���ہ�m6����9�KC����ơP��=�3�s���m�5��EϹhf�2��z/��1X��ژ�x��U$c�'�� ��VdA��L�)qJ&<@�F��Ά��6A��r��v{Y��	cʔ']c G��=�*I�����D��l\���o�?�VR˱���d�e����KETB����隞3V�_���ш�^UԒ�c�?���BUao��{9��o=���Z��: ��D���R��.w��CIuv"L;ؾ����>��3�e�4��o�l��Dd����>�p�� �t�-��%�&p�p�q֍h�"��ln�~Ƿ�O��V�:���QO|��=��Rᶔ-�lw��Hi������ݍ:b�p|y���M���㠆){����gZ�L��拺�]�Í"`�H�T�!��n����3r0��@X%��-G�8��m�j�r�%�-[xbHH�?@���G��� �o^È������kL$�����:Q/���"���zD�RvL�c�,�G�Ԕ�az��q�#��'���˃�#��(��ȥ�yC���lgԠqS#I"*le��"H�D�<��y�v"K��[�c��Iϔ���̣#��+y�k'	�{�P�c��-s��jw��.f�s���w���y�N�t�����>YW��K�ߍ�~I��SN:�� �UeA��R����_p»^(���@��KF��q��s��_�F/dð%��@���W���-橬F�(@y.F�l6z$�w���o*����X���$
K��粌�t��$,�p��t��k�x��	��u�U�I ���\�7�ӂ�4���	om9�ylQ`��P"QڶL��Y�e�ҵ�%{�yf�(��/�:b�']^�]�O�F�����N��yn�*v�*:���������s)�#���-�����{<���s�M���q��t��k�hј((7
����MU��e�N�0݋��$B�+%�÷�2|���_jE[�`���1�< ���o%J=B$��9g7|
��j,:wA���#����7�T�HT�{5Z��%^kY����ٌf������cu�����tS�w�hb��E����t|g6!���F
ڷ?K��*���fa�H��ƣ *u�����^M	zܱAHs��`���9�g$
Rg�e����UQ���e��i��`��Cf���փ���)YcvcJ�)��6������u�)�܊�n\�t�O�Q��S��NW�2G����}B�~�H)��F4X��P�P�D`^��d9H%!�nC�k��c�^b�a��Կ�pA�����3�5��#�"��/��.���zc�YEB�C�/�"����atp*ΑS�o �����b�[b
�Ј�s��
e��xʰ�B������Ń]�����a��pͳ��ע�I8}Tr1�U}I��Fo��NOɻ$�Z�:��Ԛe�2Am3�
4g��?�#X��G�3�� /�!4��p�9�l���ldvy��p�!����K���,���Ic��pfÙV$�Gٝs��vH+k�@�D�T�H���Md�xQ|���G=}��`����*OA3���a�T���4�e���g*s�w����`�kB�7�e퉠��1������2Yk��t�b���Θ���9[���JX%;�Г�\E6x�#���WdG�Ə���T	7���|��p�L��(�~����u��r|�Cx~�R�>�.d�:w���'1S'Gs#�ß�t@����~xp+���\"���V��}�"r�B��_�P�c[t��Z�Y�z\X�Yg)L��g&#�����Vͦ����Y9�_���u�1#|f����_�e���ٷ]U�e��WL�ճ|~����ms@��A7ܖ$�C�n�I���U2}��(�)�bjdŒ�ڂe1I,�̥/q��) G��w����:�N���W�S��}�O"�mEh|_8��Di1��p�U.�fϥM��L��k*��0Y_�a#x�s���X=g���'7�2*�B���&yY���//��i��Y�z����_��|��[�3߾�z�f�hd�?bcT���=�E�No����mw�"����Gˊ�H>lz^'_�M�G��j[0�Q] <
͆XȞm�_�3��|+�s	�c X�-��S�����&±kB�x���c���~���T�kY2[���l���G!4��\%�`BI��6�)�ɺ���~���T&�"T3+��"�~����Q"��l��F�i���l�#�����mi�������̻*QCMv�%�^ �b	��1���ػ���Hj�M��t&(ơG��T=b+0�����=a����>�_fF��<fM���d+#�~����?U�۠�����#�\X�E ���l�N���G�Ri��Z���ơ��{_��.zl�����\v�fY�P��,��=��R�e6����7(�C�T.�A� Ы5�3��-�2U*NQ=�<Q3�r��E�]�����޴s>�x,y����fF��KD~KӚ �=6�	�گ�(MB�4�@'��><��������'��׽n��#�x�K�l�C���>��elb!��j��W,"��\�!&�Y�@q*�R.���j�b�[b B��H 4�tJV�i�y���%��cG�;F;�,[�DA.��_��N�s���$1���%+q�aQ�:�?�/��'�{��5I�0ֽZ<�x{����V7/�⽑�B�n��74����]���h�)|� y��~�"r��
|�	Q%i|\��//��01��o�iC�"��m��gZA��}��m͗�^홷��Ȝ="a�L�!��]3��+����h΂xЉ�]�K�t�'w���!ܽ�p�#�q�t�b]p��I4�ߎ����K������)[G��!;]7肆��I	fӣk�|�DB�����o�5��0��Ȁ5���>g)}�ڤf���)�h�$�6:�=gZ@`��1Y�5=k�����GP���kS "�Z8��z*\����A*��Vk/�T�y���AW̮�})�C=�W�;v�V������� OE�Xj�Zv����e�vy��]<���q�
"|Q3v�E�vJ�\>�p��R_=�X#[��N��HJ��� �<�����*�1]Z��2�f���w:�`��ۮ>�ς���]�gڣ�!�E����֜�<�ׅ)���r�ޠU�ϒ�L�Oh���]��	���9\˿�"�H����5���a9 &���>jg��I�XZ�??�`����Hr�42l�����4��
��<N@��`u���:6���廷n:P�յ���Kzs���&�L?�3�j���4F�5���I��*��*�v6>k���5�X�)���۵N:��3��<`�+��D�����l��|\�dcp�#w;=o��7b��B�Ѓ�K�~���L�3�mZ*�]��^�}OA���F ww�P�y��"Gf9���u �i���
��[i�>n�R�$�-���mȓ�9�9E��UC��W��k/"��	
�J�aY{+�Ƒ���9q�`���i̗A�I��e���z-	��f��O�[4��\��˿k�2������}�әm����?�89G,��
A�Q��+���h	�=n$�p0抝~�����d廓�L��׍�f�.C�-�[퓷���yJ۵#/�g����"���,���ݲB0R� �jfFq�� T;/�f*��ذ�N�e��!2���ޣ�$�ۆ�(����͢%�ǈ�8"P��w�x�� �'Ifq=�`����B��� �c�y�)����*��n3b� 3�Lv�ur�]�٨����@>�*�Y��B�黄9�ɜiGuO��n��	Ã��yJeq(^������BOY���֦���K� �`��"l,�g'"y�$����	���S�8̦�v�zƨƤ��	�H囆ߦ�(*3&�X��u�m*�}>}jNW�W����J?�Юrm���}v �8Z��
^ԍ�9Zn0Be��#f�ZhC�hxNy��a˟�fؘ���5��j��c-��p"I��n�	!z�6p�E*?ad釴 ����g/�+_
�,�����4�B�3t#��@i����K`rVK�?a�]�n)Lˁ%��"�nӊ+�� ���o���ҥ�:2��U:������&;T	��)s����_�����]�a�Q<h���Ȅ��U�_ĭ�ϻ�M��d���P����&B�kP*{d�rʔ�_a�By��ٝ
�$V-<P�^y��<9<�r�? O�R���;���\���~�|PP�B$F"�8�/��=,��L*�a��e�%���J&Fz4a�� &f;�|ߝ��@�Ta�o$L>t�J?�xS7~��:U�I�1�R�0)��"�GP���},z��Q�]mP5�W[������A�t[�^P+��mjr��-`�Y`/�r���%�Q�Ui�s+��ƹ��c7#�L��S��/�1���R�,h��c����v��K7栔�\��"��ڣqAj�v�}\�.Z��3Q��ƛ=$��!iL;7� /�������h��R�B���98S?�F7�g�f}�p������[C����f�Ά�y�Nt�&�27w����v~Jqu� Mpu-T
(\@5s��P���	*s����,�=e�����F�>�=ҝ�_����>8^V���4'����\&v����8�9O9�� �m���Q���1l�'>�C���m��E��D���&-��qM��W{.�3��J��N�'��
�H������P�\�3�]��ˎ�]-�Y�~�d�D�٧��:���]��|݅���r�m��w9S���L��qќ��0��!+����^�F?҅�X&�%�aڑ����AY�Zj�"2>�&��kD^��i���4�!&"uu�G�p�%D���t{�-����0;�;j���Ppv�P��r���u޺LNc��b��� G�<]�����_G�yE9!�����m���y����zDm�Qg[}��	��A٥P��(�ي�7� WN��|
����=���ZL��G�c�B�z������&��0��E84��&=G�&]�g1?�p���4���l�)�迣vf�Ŏ�R�K��'���?PbK��$6s�D'B,t=���<*�ª7��r��#ԫ��g����om��g�Q��y�qc��Yu꼣��o+ �����F�n��O�qa�?���Q�O��w+���D���%�dXٮc� QJ����2��OD�HA�ƀz�\�N

E�tc(�I�O�&RZa���h?~Ԯ�X,�D��೓�/���T���/$쇴aAk����W� Gk۟����/��_���	>KN��l$�	�::�ʪM%�j؃!{�K}Zß���5r����i3�G�2V�zlk��Q����l���M�p`H��D�R�a2̀n۲�ږ��"��y��m˰d�3�|m���z���Xճ�ŉ�
�YpAI~!1��ϲp��'�Tv����xs&�6i�4�m�ePY���m��$z��H�$��n%��P/v��t�����$�M�K�wv:��\,W<��q
R<6���K��i5��U� 4$�PV�o,a?I������":}{�l�H��k�7��+ŋeT=d��)���rn�KQf�c ���z�r����ǚ$�ڦ��у����#*���#L�j�$��z\�L)i|�!=����ʒ�'w�����/�y�WkM1�t'R8m��t���.>ﰘ��ij����4-q�
� P���S�NaJI~#��oŋ�Qׇ�Q*���h��p�]Jvb�BD�(���?%ci�v�צ�Mc���)r�Z�LK(�<y��"�=���4��T2\�|��6���j�\;�7�[�%@$_=�o���p;��7oZ	�+���j��a@Ӱmnv�ظX&S���9���1���2�ٕ����e�Z��J2�ꭉ(�9�Ր$~�a�"l�LK^ŝ1��7%,�Vծ���U�A�,���}A��'<;,��.&�ףT��T�05��riB蜴|S[�H��G2��N���D����|��la�#���@k�&�i�SQ�@r��UB��v"�	�=��vʱB�����Ӫ�O>�p�MM^�F�Y\,@u[ca�!s�?�D��I��B����m4���Y���?zĬ�4]��+J'�v�7fz��n�ԙ%�d�F5��ez��q��r�fY�ŷ갉���:0���
#��\�caN��Z�%�k��\{���Se��Hռ�ң�le��0l�K�Q����Dͬ���c�ڸ?���S�&da׈��;�^k�.!*�Ŀ�Aa���~:o�3`�(3�+�9$�����Y�_��8�.	���6���� Ai��&1��g���p����:F�l���S4�E�'�@P@�e�ce��$�6�rY0$hW�������a
�4H � 7X苩}5�@h��g.4@C�	�vR,.�� ~���|Zң�N�il��%�8��|�o��8X!s�vnR�{I���έn[�.M�(&�d�̠���Y/��t�ɓ��t~$ˮ����La�Ȧ:�-N���e��'i!��o�8oٜ�]W3��h?���U��}�ѻX�9�hJ)[�m�{9Q��on����	�W֮�1'��ú1��R7��7�xzvo�k@˧�.NK��f8-�h?k�6�G���LQ	��Ci�d)���ߘ%��
�G��+&�=c�)���h:��na�[F<_�e����v=ȏ��bۓw�_^[�Ւio�>��y�Dxm�N�0�!�r|�e�q��⁁�'����&GN���`V��Sl+J�]:�(��ǂP���؇�	l��F��)�	Nu��A�L���%��L���3�JPq6,(�"��~<�Vε������.�Z
@yFE�-��k��B����ﴢ���e���M\�&�R=d�WB$�8*��[�A7�f�ŮDeRo�)4�
=k* [m�]�����k�V����y��qm��G�Ic(d�;~-q24׌8����f�!ߜ���<`q��o�&b����T��,� Z?�I	��f�n��q�u��|�P��C�c�͕Ck�$$�Y�5��;�d�%�=���ںUob$��������PNS+w��,���Cv,�q���?,��d:�) �%f��������õ.�G|�kAp]����CU�v����78$�كp�2�ƅ��\��YU\0%A3��o�^��8��r�L�~��}<S���l��|Ҏj�8�'	MY�a��#;�!\��bZdX+/��b���I{Xs�%��R�RlNV�QJ�^��)��HF5��o_���J��׸�H�������j�u���A��i�,����CM�MBI��:^��5" ������� �y�M(����(���D��j�-8F	��Q��lP���S��� ׬�ډN�Yߚe���{�����{��6���r$;ʥ���ӧH���HMT"2n&L1@@#G� �?Ŧ��'���
�{�xaþ��;����D�v���'�#��M���n@���A(^d�{	+f�J�a�]�Br�B8"�A�K��۟�S&x(��I#0K��Y8Mq?�ŧf��d��q,�:�\�/��c���c�Z�2��c�"��������N��m�D�OG�	��$�@���ٹ$ � D�f��Ha���.�;%��J_	!�KY&��Dga�`Tq��>�8�3�K�3���\���Q��ֹ�:u��|�tH�[��z% o���dΥJ�L,��J]K=3��L#/�O��\3�j$�u&)<����lZ2)߿��\�T���ی�E���;�'�U:��G��L�l���R�m1�`�Ͻ��O�tN�`�v a,��;lL�HH����b�3�|���<�Q��<"��Yc�I,���V>e֡�;J�W��82/�s���m$9�K����f��Q�2�9I���+]�i�r������
{L��R��������u*-���J�&���@���B�R�X&�£�ZNj��Lm�U����<�||�MBnʟ�ڀ�1B_�4��ӛIa��2l�����������bx��Hk۠@�1�|�T[z��
�h�?�1�bY�V�`���Z�(?{@Ys~�
�쾗�.�YAԂB�I*��B�i���DT��Hk�Z#"r�0AE�f
M�N�h��Q<�+G�GM/5kJ�v���˪E�	.��fq��� �K;r���g�-7��H��wi��V�^ ������R�1cc�P�ܜ�H�쏶y��ht�d��ZNi�d
�qt:�>*u�K�n�Yr��?����`��;��=��?�{yz�"�������[%�'n7EQ�&y���C�e���P5Bg�z���Ȏ�wP'[:���1���f/O{<HXg0���ܜ	@Ų��I���8�c�S��7x�g��r�ls�I����z9Li�R�=f���3��i����y����'��p�^e'�b+X����{����o<�y�Ď�+��.d��/̺l~S^n���ԒK�Kt�Y��O�r����n��̗�`8s�l��<��F2�r��#����j �!v����&v���K�����GC^�5�0��A@���k@Bo���=����x1�(�	j�8_;��t����M7��O�&�'\����d�*���Ann (<�d�O�ս�X\7�@��۳um����(�wN��g�J2	�x�@)ޣJXZɊ�b�7wAA��D��Fa��T�җ�*j��]XV����A�iԶ�3����l�V����6��y�g�?��L������;	�)>Wλ$�M�]7a�A�f˓�r���6�$7�$b�Q��oc��f���u��TI��)]N����<�8���A�D�j�rDu�u�S���:Ev�nt
��G��˩���8���V�"�7�m�KI]�k�H�L��=������������VI���}Γ�ʭ�.ǳG����U@�A�	�N��V
��㧀G��^�k����a������guc�!�P~Gq�L��tiU ��G�؀� :��4\�#]K�΃>��B������*�j�v�������%��\)e���2I�,!�EN����U�@�#�х.P��v�@P4H
>�~���S<�s���.��r~���~]����� U�+dhF��������z)�a8�D�~�-,��}[��B�K���r���w�H9��Q�&��Q��3�]_��cS��Q����{��b�ȕ'��R1pR_�����\��w��1@z����U>Q��HJ~��"o�k�_�L�v��6,�z;{��7o�Lģў��o���AMzM��;L�5�����8(X�{�#�(-����ȍ���f�l���0�|��������_��**�]��AIr� �'��TW)�>���C�^��`0��T�ܭ�)bqY{�^�Z����<d|��
�)�ڭ&@P��w8��&���I(�|�M����u@����D�L��F����i#��t���O<2��F����E=L_v�Bm8��"��Rՠk�e�UH�����N5��ˈ=��΁��ϡb�.w�
�K�/�Bc��]+��l)dv;�T+r�E@����T��MI8�U�$�G��e�-c��X�]�ߒ��σE1��΅�y���rT���<��$��
�q̤�������ޠJ�(�W<��������s�<��s�U~�K����!�|}ٮ�=���c���0�q|ܸ7

ՙ�*�&pC�7Y��}���Lm,x�pWA�a��ߴW>Y�*�v�c�gjD�n=��9���1�Fb�ຯ�Ȣ<�Y��괲�`��*�||��7�w�x�F6��3'�M;wP�8�Eky#�Jh����0_�V-)DP�KK�N��Oo)��L���I*܁~(f@��y��y�P��R6[�&J���M֚#0����t�da#�^���a%_��<F�m�~Ư��׻t�E&Z��x�Q��_f�� I�Uc&)�c :d ������K[̨(T�����7L��6C����Tg8��;�C��o9�T`��ƾ9�{o�6�ǟ�;˒~�����v��ǒH+P�	���E��;+翑ol���0�����nRE�
������lg�,v��J�A���#�O�V쫤��4�����4�2��h�4m7�4�o�l�����`_�@���*'��4��A��`_���9{>=Ja���d>|v�OC3��Xrd���տI
qӐ�:9��:��b�()�f"!�$��G3�+��%V�I�ȅ�],��J��[�ю%�<H�<�� ����We�+<��k�E�!�8r���c�0���YU�S+�V�/�w�Z�Y���CF���#D����W>�)A�ֽ�n��p�1�r/����ǫN���xʣ2�$�p5qlW�^X��]�h�PaS��k|3�L��>B̰Rd�T���PR�T_:�x��5��7����ZX���g�JG� .�;͊z�m�~����>g�<�/vBn�ؕ��q
�,L�\������g�d�|{_�ɻ�R~�=|�;��~ʨ��k�&�$�NgXr��bW)�R�O CV�+ޮsxĩ����^}�-��iJ�m���5��SNG�E�TN<�.�^u������xѮӝ���u	�P�֭����
Y��]CY�Ǻj8��_�.�b3��s'W�D� ���uL���|�J��P���p-ٳ��D�� '�QU��f��&�X���y��G9q�'1�	���(S[��UU���w���.Pp}~�6�M�{fI>�g�����}i�:m�˛�B��T.8Y���ef��0[?���o���ܐ��WoQ�������+%5�ye�} �+�L�DU�o�%gc��PM�Ab�kʓ��HG�P��dK~L�t�5�כ
�]`h�����Z�P���o���q�6@�9d%U�t��y��39�3���S��e�}]pen#5oX��Lx��R�c�!#q:#���2"�l�b�����ţ��2�=��MQʹ����^9��� �bA�-<A!R焫��Y5O������eY��#��5��~S{/8��C��{g�8]_A&����'���f���*�n�.�q�d��..!�{Z��&d�e^J,q�E�NlV��`�; ��\#-������f4�����R��6�d{b�,I�ˇ1ݣ�Gdb���������S�-���T����Y]�ַ��[�w@&��*�!��g`�ף�r}^�C���M��62�+(�J~
�[��b�;?�T�ւe���HK�o�����0�k
G'=�+�����[,�^o8��T+i֡�n��i�j�TS,��������9 	Uc�*�j��)���K�!Q+;�nsN:��� ��i9A�0�&��Z;6���ь�������W��k��n��XJ�^'����š)a���>IQ�5��)�E�y���o�N�W��[3��L�j��2I!���_��x�8��]�8��*��n�q��2x� �����z:�Zp���w���#���_{�?K��g��9+�N�2��0/�����9��^q$�S89��|��Vێ=��t��@u�ҷ-l���g5�Np�ZSƺ�#(_���������	)�̍B�#��;�c�u�D��..ԉ�0�5�*��[Rg�<��F��$K꺞�~_[��6�o��%!K7=�,3�q\=X"��up2y��8�̂�f�/21�7��s�Lk�$����z��NO�'�ݒc�oyR��zT@]�!ꈉT_�B�,Q�$p7c�_H�y;tM�-�ٶC�Y(�T<�_@3��VSX܏(�J'/�t����c�6R\���:�$�B\�� �>;�VT'65�:��v=BK�H^K�;a�-�����-��O��r�׶�%�����s�ϸxd�}2B=2��]��:�m!'���ՙ�c�q#�Cm)9�G���2753���,��i�s���ʀ[�%?�j���K΀t��W�ު0(*ᚤs��o�ӃL|@U:Ee�/ǄK�������0��Y�;��L�v�zESoIښrBt�p�+�ة�|>�?壇NQ�\�Iy&I�s�]Hő��/Jw$����h��]oXګ��-�������߻L΄˼JN?�.M����fVg���8�%��D��(^�7Tp���*H]*hf�";�6`�}ZNS
;9t�T�],+�T��g�+�|�k� �KT�FY����C��<W�3���%	����8dS�s����E=n��g�9���5�m��s��b�K��TN��ߵ^��P!�,5�U5Q^^(��܂�6���ߥ�!b��Zc��.���Յ�#�M�p���q�1y6@�q��"��h�x�~�w�Y\y6������摭�!����"��#J{�W�πC�� >����yYe1�W�R0ɩp��h��	��2 �M�E����|e<»+N�n4�T�P^�������\)hZ��6��+�ӿ�h��\Ȏ�@	r�jds�V��Qj�/���H7�gP���*�������@�6$U�����qr*�t��
���B-$����D`SH��°Ә�⮾��}tR㳷�,Q����o!2CdM0Ӳd�%�NY)�'Y�T����ø�9�	���JoϽ�
ʹ��5���"����Pa�P3��f- Ha�L����p�#�#�5#t�)E��q��`;�A��(V�c�֏�@��nȩ�Y\꾈CJl��)�0���lC^�8�9U�a��6��Wҵ?ʛ&Qz�)x�Sl�)�UV���1S�KW!��X�,�Vd�H�,ulӛS�'�t����t���)IX[�_[@s��bZ�w+��b+*���%Z.+�1$;���4����k���\ʗ��-	�E�U#F��B��!4S�0_���n�KS��E�v���⮁u�n�,��#|��ڰ�]�?h>KjYFR;�a�U��ADA�T���^w�"&�����٫L��N( �k)�%1Qǥ�$�9]r�EIY5��᳧���$ �{���g0\=;�&��K��`\5Q �=��s�qbޮ�j&�Qㄩ)n �/w��Nj��0hN|�W����2w���n��K�Ŋx��ĕ�Ρ�ۜ"�s�JՃ������λv���� ���hه�C�_��T�+�Z��w������sT26,�=�YZ ��Y?�7		)��Xar
@���v��ڊ�1vR���1>��Q8h��T)k��[I5
&V�֤&�Z�p�Ц݉�.��_��� ������<兝Z�gŁ��!{�Gxұ�Z-4���[ ӛ�!��}�'	���SՂ�b�Jt��}�R�(���?w�A@J�Z	��͆��c��H��Z~�n1�uX/���(�d���m��T��ۧW��k��d:hۋ��`�U�C�`�0�����6Vޫ�_����N����!�e*�5]f Hw#�_��ɴli��o�o�C��g������g?��#]&���<�l'lř�b�E�=����y���r~jE�i�c*)r��.���m@��:_c�����No?�T���zC��󽓣{Z���}�4���v^�Ŋw�b�?Xgΐ�/���JlFZ�D..��Osy��W��@?���~����$��)\�Λ��ҝ�X��"
���3�"�o^�l&���<�.�S�_��R˓����щ F
���8���-ZE��u��O�֒p���c��A���'3n���U�h'T�����nQ���a�a�
~��OS��掿^B9���i^[�U,0��5�7ö}v����M�cȆ�U���5C&��bz:���P7.�$b���IF]^G>��I�wn(F �^��Ցk`+����_}��ʸ����?/�� �+Ka�CP��h�i7u757�p���C�bor��K�ּ�	��^���������]�j(K6��e:G�x�����2qx�dp�*���a�J�Z<��D$D���;Ͼ������j#�2�*�2��CR_*�KM�V���c�f� ���a�ȍ��Q�y}��F���zŜFS�v���g�ġ8e\���7�um�;��x����Q��-{��j����K�yP�aL��HZ�n�%}���WN����ⵒ�5E��ɱg�$&PY�pKQ�k$�i�b���z`�LSX���ߤ$���o3d.�\*Rx�˫��
~8����s�z�%$��ԛ2Qe��WjcBc��w�#2�G+���]X��hz�y��<Mu� 2��Vy��⤧���}������ynfr�h�cU?Ё����>��GO�'[V�l�)T�+��C�w#"���I;6v�P�1�'�
(���j�a����"%� `�G��,g�L �jD���U��bݮmdť�	�S�]��L�9�`e�dU�g�o#�p0�՗W��X��!|D����(|8�S���$X��ض�%ͧ|�	�SOR��Zf9��>{^�ܰvy8�G�҄ F���f*ĩ� 3�Dl�lP!�/Ո�/��=΅��4V�*Z��׃�={����[��\9�f�7fbg���*���:;ƾ�^]�ۧs�����s�ܢm���JI�S(=���n;��϶���!�ȵ��":/�i~�|0�������CZ `_a�V	ӿ�8�m>����ᭉ0p���rΠ1I�d�ELwN�����+@�O����U�țjN�\ۏd�$Fg
R��J�XC?��%���9X+~���/��_8��F�L����.�\�Jj˝�&�u˰C�?;d1�����QL��x�F��š?{/:�m��ܶ}���ѝ4z�*��G%.1���.��{�����Vs���d�J�ôY�a#�'Ɵ��<��lqŲ� b����r��h;3���i��2�h��N:��}��5\���܄�;�q�j�LA4�U��!�U9���M��dfF3.?��w�=��$����V�7�Y�ʼ�4iԐicYp,�o���5Q�L<,/�����Ȃ޺��*]���c>H�����]��������ئ|��K����f&Ⳣ��^pF+k]�/ND���Jt��U	����A��1@�����p:X"�^�+ޝ��k�Q�qh��Zg"d���1y�;Б�f q���}A�08b�+f��Ԧ�)�}�dϵOO��+"�9w\ȱ��?6S}2(|��ԴE[
�+Ɍ(�Tͫ��.ϖ`��5:Qh��+@�����m�S����#�$���d�� {�C��4�Gl�g���"ySm��M�y1��� 9 ���]�y�7��J�;?3��Y0+�\��2 h
á�F�w8{�Y����4��������T$��-T�0k�+��K��p��;�.zD���-�����j%�	n#�g�J�k�A��l���٪�������M�T���B�rxIA5�d��00�α���5?���9��lAq�(,��K@E� ���(���ұ��w��n�*:kF����� ��F������G����d.Y6��Hq=@s0��p�)3�&��˒�w��.\�t�N�Ӵ{)pݩSG�5l!=E���8
;��������� ���μ�}���.�)Z&��QEIX[�V!�n�>|W�w@<C6*o�i��9�����Q+6�c!�m#W1��&��X��*�AY� ��e?�#V�3Q`~\���~�$�S�bZ^'v��:�u��(m�:h%����ml����d�c����?����FP�iv�h�Ɲg��K���-�C�7(=+Pp�+���m]�=�%��;���S�fx%�s�����ڢ:���2�O��IF7��n�&�g��{�s��p5��X�y�i�羠���ՠ!ᭇ<��+��
l�XGu�>&���n�U3��`f�m�8���𞶜�D�[_*�1/����׿�?��Thը�4��G�;9 ���e�³~�@��ɸ/M��k*Y.#�|:��W��.���z|�ސ���������6{"7�1���+A��F1mO�V-9�Hv����6'1p,���`��eYχ�M
ӽ�c�f����o)��%i����@�ܮ�UT^JKԛ�9>�~P�7//�,U<8I%8�h+��1��
{��S�j��V���L�^0cY�Q}�BU�U��z[3-56G�ؿ�r�(�l��:!*��񳂎ns�7-�!a$�m�V�C�φb���'�G��/1��:�H_�7K�w��;Y-�T�M'I�ؖvyb���mC�ޮ�dQViy�/�Ѽ�� �#�����NW2ʦj���;O�S��a�Lx��oU��v(-���A�u����_L���u�q�H&��(�y�i>��J�MY8�D�&��^6���w$;!_���%���b�m���G�Ի᷃NIR������ܦ#��Ry��$��7���oҶ����9�j���ޑ�#�<��s"��q�^FK��+д���mO�=�%A6X57 ���9	�Ɖ�c���+���ؙ�ҙ��M����\5�;Vv�X�V�<bg��D��ݜ�M,��AGl�Y,����e��-����՗��f��G����+l��� �RD�\Jf�fi�z��^$�P�h'�v2 �@�+����+ꁔ��w���ƫg��"\\�%՟+5���n8�"ٙ�V@rGMW4��N�_��y�RwOF��D�cߠ��َNސv�}�Q��o]��[5"Z�hyM�<9�l��.�L�<AZg�f�"˂a\��c�@���.����̲'�&�Hr��7��ǉ*�=���)Z؜��A��CO�=�v=3�Z�ZQ��c&�9(�Db>�x�����|}������4�X�{H(���U8�Z'h�NzB�	�a���nmu� ��M��ڱ�_=͢cuח��D$x���LV~
�)�ү�tJ'*���d5�ƶ�AT!F���m������'�.)��ڬ���	Ѥ��@Pǹ�,	̷]ϳ�jm����*�M�tR�Ѵ�:��;)���lrv�T�#TH�خ�B�1���0��+(,�7z_������$%I�k�f�4�)�4���M�!��w~���u�զ|zp���v	ks���ڄs�:,Wxi������}�BO��I���B/\��h��� ��s~��Y
+���
Ŧ��^I�r�X�?�С��J�I��nޙ��*xI4O~�}j�����O Ƨ�E���3a�����6
��D+��KR��6��1�>�,k<�c\��!K�/�"�Β�y,
��(9��U{H��nBH��G�v�/��R�L㊔��FS��`,����&�ڷ�ч���|����=�T��G������<�5\"6��Wxao�4pP2�����1�]H�E:��s3��^lp�R�ҹ�`�b7���HtU>��&���ĩiو�d¢�]J���"�a�cWP�d���P� ��sJͲN�ax�ra:����=%Y
�9S=Eh�)�␄�fm-�vij��<T4��?��2���Q�d"r��	 ޱ�}<��'���Y���&��_�{h�əA�Lf��;�><��,�Ux�9&@�e���#i�j�U��D�l��(��˺Vͻ���	���* FJd���͛�$��rw�d���j�c8�5z@���CћCy����$1wx�u���e��o[��a�"qQ��|O�� J4�\�u��|Q�b	l�\�H��j�u�a�'�'o�e����dC ��d�BÁ��:�p�������r�@eVsY�q������R��cݨ ?��oz�#+]=1Cj��wO��Ї�/�H�W%��T�L/40�ç�(z#D��͕��g����5)�N�	ķ���,�����n�&�<r��%v�H��S���I��L".E�s1�l�E�#Z�~��e||ŻA޶�0r�Ā�e�����:�2���,��nC�Tq�1T����HY��o���ܜcaս/U���Ĥ�
���*;1�ڢ<C
��f�7)h0��rQ��fm�0.,S%a�i�+֪h����tCQG2q�􈨴�HJ��ҷ�4B��$�FE�~^@3���������曑_~`[���(�u���������mMo��<��ǥSH�mX�_��A;�F��K��o?A�8�Jf��X*�>���P������՝9��������_Td�b�')mI0�cD���]����F��y�f\:�)<���uT�`�c2S���@����*�+�2��lYv����r���oД ��>ɻJ>��ĨK�d�^1��m���4��E����0�(��|�7VÕa�d}C;�c�C.���0{,֋a�(
��e���Y���^CqsV��.ʿfnp�{d�˦�j���ʶ��p�g���)m���a�����Е�v*�-�Qy�K��E���q ��nIT<�4�!�n�j��c�nd�C��/�4�����f�(�@����m(�!uCN_O!�|�Ţ�%c����n,\�EK1Awf(>T8}�+B!�؊���O�#^<_�6�1�y�T�_dh�p�n�l�=���l�����N�D(\��gZ��K=J���j� ֻ��>W�tkj2r~��10޸в��;uCDǷ��
����0ᑿ2+y�̊�b`��B�����9'�+͈�kNq�ǧ8t����qc���
RJ\�0�O�6B��N����!�x=ĕ�7��Vf���!3'�Y����OH�1���R1��)CkЕ^D{�>Nם��͓[��Ue����-��<�^��/}VzY�O��^
����QBf�A�eK�ݷ!�l𧹪�,D����K-,��	XM]I0�Nu��aZ�� Otg8� '��(�����,0tV'��6][�b9���SV�F�,�~�g��2g���X΃VPu��* ��h�l�=�k�c�R�֜�4,�|x�W|�n�@����y�?����i[q�S�f���$;*�>4}�}Y��X^�Ë$�y�C�Z!�ml�Tv�!�7mǼ1N���Trm]�?S�4��q���k|r ��I�U���Czb:n�����t��߇���x=\(|��DMb�8]�co�]�Q_���Ax�Q�Z������,��.��4X�ԓ66�c���=�<�g�ݰ����~P)׶>&z����A����u����O�]��������~��Ie�\�?o��=�P�:�y ��+&=����+{r-�_�s�o[���$ ���R!����t��L�o�}�-�I�8��q=��rCAr���ͪ�h�|/��v٣�M�L�e���>6'iqU2����Ռ�../S��=���"ZE���D\ �\�?ݚ��j�^��:i����R��6+�;]���+R�p�SJ֌�HV�������E__w�[�O����d��m}�_�i�H��XqZhŹ��Y�v\r*d���w�K�u�;�"_ƍ�}�U�j�����=<JZRÙ���"�B.�e�~�ۦM���!=���ٌ��q�;}u}�W���_q,+��$
�Ag���֡�$��h�/��L\�#[�[k�/���ju=��l4��&�~m�v<����HX��A�H`���9jr�@ĭ���J�G��19b�P������o���)�'?i��e�;��)�������t�7g�m�b]	��%q��CC;C`�1�}�h-��F�\G��!\��z��GC�����0[�L�y<\!�l�2���<v�ش$M�#s����@�o���s{�i�}V�?B��I�d��=&��d�Z(T�X���~i >�)D�0����D��+J4\��MnT]U5������%Q�j8,�J���u�4Ԕ9�{݀��*�1dHsR�J9g��
�Xn/�㯨��dKCgw.��8h"��Aakόy�ϯ��7Ȝ�*/Q,]M�����~15ܲ�W/b�����=����wyxvԜԇ���u��V��8���O�G�����$Ar�搽l�A�/��qk�_�9�[�F�0�r5�����M�/~y9[��hK���<YWT;@Dw1�^�_�>��^&"�k����~W��S�` ��W4����DT(L��i���7�5��·8ԃp�Ǒ�=Q--(|��@���U����=~��.;�.W��3z+���ne?�쳝�2��O��o;�"kǚ['Z���d��]^O�8c��PB�N2f���b-�i.ϗ*;z�~%�6��$��:�s�D�h��Y��M(*���p�lv�v�0�bV�7f�ĉ>�q�w���#�D&32Z��"�B���
9�m�ˉ������[_4sW�V\z)7=��ȇ����(�jd8.6��5������09��
5 `'�3�z,nwdd�sWK��=S���V��m�n8}�=�WB����!��&b�0�����x�
�C}��&�Rk�Y�1#L�O�H1z�أ�N���}c��!J%�A�8�V�Mc�U x76/`.�ٖ��������Qi��f���P�v��F�5!e�5/4QAB�7O�|y��ĵ�w
�Co��?��ft�����(��Tc~zdЦ�j�'���]޲k@<�]�B��d�vKCQuh��ً#��5}�-������F(��`]��Ĺ���2�zD�g��z����S�n$*u�!�
s�*3�抧)�y�%-`��s�~���R]�f�i�k�%���+�	�����U��t�`<+�/P1=>�����ZG��9+L�g�(�����,ewR�Gfg^��`.�&��D��N+�Q�k�Xc����|R��Xg,�2.Q�_4K��ޭ/�FPqB.d@ZY��^D�S����i#>s�ZJ����f���:�;��g�xf٪6���Z-%���&��,L��ҩ¼�x]��Q�g��U�S��c��]�l�Uѓ�ߞ=�4M�B��j�l;7�˂C��u~��)@o�?���ʳ�^�KhjT���]xޅ$r?�#G:ӴK:_-�O�yF��
J�V��5��dmnD~��3��F��Ϫ
Zi
wI�EP��� �r��f���R {�2�7Ndz"��2���:o<y}��CX�oq&��L�#Ƿ'85����3�0�L �R����%���I�Z�#���+��0xgT=�J�`��_ [���" ��h	��Kk���ɬ��F��@�i��Q����BƵBTsnQB��E��@<ѠU����B�_��ؘ`�p0p K�>�ܴ���a���)R���C� ;�,�0���̓�XEAnTJ����oOc��;� w�(C~��LV*ic��Fd[|R}X("�AjO���ŊC$)~�Em�bL��o���tn��A/��i ����:,����?N��+v��e{��ez�sd��ҊW^0[1�e-XX�6;�I���a}a��>��m���\@�4xu��6d��e�m{�gd�_aK��`i�%X����J��y��m���@��5d�(���߿���<y�U�D�
h�]�kvޯ���y˚�h��C��EP��h�mJ@�
�xǣ���/eR�<U\�AT�|C�	�0 �mOX�s��#! yk#�>��|�m�&~��V�g|j)MY
KhwZ�*@�)�uT�L��ǳ��y�g��4���O� ���L P�a��ǜ7�n��:(
���
�+Ɍ�9;V������.=+�oC`��qnJ?Z�sq;�8�oʝ٢�'�A�O��������V4hk�_?��dFD�w{=��V h��i!�$l�i����r�J?�Ց��j3Qm��0Gu˾?�&�J)�?��]�STқbpw���|�f]2K��cH�P_w�04��퓌��+C}�B��t����=a��A��ѧ����"�{�Y>]�%���Y܎�*ݥQ��[�\�A�d��(�CF���C�h�湿�E9��͟}8�o���X+NS�>vƹ������ �	D���Y��QHA���T�1u���F�	�sn��� Ţ��S�t|�J�p�/���'�{�)nc&k��Q��0��J((%��e+�*C�<�/ƫթT�MB� �`�6>f&.SD����+;ӑxt:�.�ڷqt����+�sj��gf���A��U��6�6s���)!a�u&��3�N��#�&���Z]����+:\3�Ć��ezą6��'�V,��g]}Q��z��}9�=�#���}�\�E��pG6�v;�� ��`{9�C�Y����t�t"���)�"��w-����2`� `#�<@?+ͷ���'�&I�ء��f.�w���яi���3����kH<Z	�rE�'�EԈ��}rW�{d�>N=˻w��$z��5��t�&y5�:J�x�sC}�O��8`C��P�Y�N�S`m�Tn���곛� �8���u�6̾z"�',��/�kҷ>Zȑ[�yu	�2Q�@�̃���K��������E����p�4��τ���d�}~X��5B�0ԫ2��⪁r^���vC�L�V�}Z5��F&`�
:I�h���l���-l�����eQ�$�_�u����p�2�B/t@�\_:!�l�v ŗ�Z�`~�����w21|�,���X��_Y�d�M7e���b�:@J\u�A�0�o��}$+kflҹsk��M"���-�NG	^����.nrHdh���4��a9w�ޘ՞ަ��
Qm�V��ka���&#0gw	#L��Bɿ�:]��z7�.H�;1t��-?֬:&^�]h������`6q��\�N��g�֫]I�3e��i�._�����
d�,�7�|�_Ew�q�Ն��Y4��"�Y?���E}�S�R$Xŀ;f�	�~�K�ą�9�WLH>��e�.:B��b����d�}���1ll���aZ�M����4{-Y�	{���)n��Κ� ��W�ޢ���H�r��U��GJ1@�h0W��Xӭ��b�Aх@�j�_���3_���F�>�G����fi"CQ*Q<���O�w.���tDD��6�G!4@gR�e3AC#����]/ �����,Φ��1��V{x�YJ���y5�5t1[��<�Lb�<n��@�����y1�[����<d	������E-�*w����|����C�s�<N7b�|�PK������C��,�I80A�ĕ?�8
���RX�n'�m��	��埳��f�����D��Qڞ��ݕ�r[:n��0N�Ug`�)6V]wN�� Q(d�弜]\��?d��v��N!�����V@��7�p���u1����`H��	�I#.Z�tl���dr��?I�R3w�'GN�.ͪ�%�~5a�!��k��/F�+|����PKC,a�p�ڈM/�g=�ü�ΥueI�qG��+
5��Z.�=?�l���a�'�.��`{�%w%s�q���v�utS��|H �!+�p�wf�Z�&�텮uIJ�h��1z�o	�\�D z1n�Y��6�5�2��$}��)un`7(Jc��.��A�*�r�aJ{-����� �De��{�|b��`n`���Mm�5}tp�[y�h�� �zo$i��Xj��Kt�!�
ޤ]��(���?ݟ^�`:��A7���X̹\�\�ޓbń� #�!�vWj�(��4�Le �e|*ǻ�͚����Zd���Oɞ+�}*U�F��\�1��ȏ�r�#B���E�B$��(cN#����P�B��RqO�7U�`���h}��M�6Wg�QI��mL�����`��W�ߟ���%�QF�-�L%�Dy`	u���0߽Y��&��ؚ+��ZqO����L��N�=�x͞{�����!�νpT��4�d_SJ��(��H�����?�.iS0���
�	g��������>�[Α�%��2�R����S�oM�Ѫ�����Ș;�SO%�a���0i4集D���q���s�AWU�;2�e"NIO��c$��l����;$^�Pf�"��s��S��K�z;Y0��������D�}/����⠇�B����x~��]��r8$�}�d�0�q�IW r����_�T��o{��͘�=��v�A�`a����$�E��GNtvS޳
�1B�v�<��cQ�Ǌ{�D��gN��=j|��,Ĳeh�I���5�3�a�<o�?�N���6�}e�p��U�]��$0kɨ�*	���K�����)�C�*u��<�ӊZ����jNѥ�?xڹ��
�,��7V4�g��`�&����B��}��m�4W�ۓ�@Ah����>�S��"��l��	��0�.�>���.�9�wY�tg���Y���6<L����� 94;��X9����ʣ���,z�Ӄ��W����$k,�r,(�N��/�I��3N>z��q�p,�eA� !_�i	Q�M������^XK �XX��PS{���Yq��@�f�(�pg��x�U)=%@�|g�b ���'wUv�ў>?.��y���ד�X�.H:ng�����k����ˈU9J��v�|m�P�JϿ�'K���c�-=����"���� 6�o�����PX�Lk���e����e!�����P��W3
'M:=E%CS���}"-�ɼ�gXL�6��"H��B_	�����B�W���׍{]��
~
�D��c��h#���]�6��z�*�FT�VD��ۙe�C��)�q��n}�e���mO*3�G ��7@�Bae��n��V��j�[`Zc�Z�Rl9Ǌ�ͥT����zw]-/v���:��竰���L�l��z�ALW�W\�~b�Ě1�ZES������D����(߻QL�(a�P�~�n�&{%��ꯇ!@�C��F���A�O׹��V��I����Z1��{:Z���5�ﬠ����	��1(��^�j�3�KD�C~4@	�����?��ݴ�o1�j�+�(�/>>8\S�����M��p�>3o�"2Z3�xB�����F4��Ü�=s�v�\������JP�R�����:u��@"�����7���9��^��m��tC�b%�pǛ�����1��Ӷ����*�uL���Y2LP5U���3�zǃ�#����yל��#p�����z�Ӡ�rς��[��jh�g(�#��Ҝ�W;Y����A[�mn3��̝í�b-�5�v��m�B:��W"uyUk�p�q��|N��Ê�[�N��T��K�H���3�>�۶b��i8�'_���d��YmPny���1<]�D�D��j�-��U
M�8'�:���q(���95���P(ּ���я�ra���}� �"f� 	z*X_w�/��K��c1�ƹ�����K��r@�f���i������z_Bc�k�k�f�{v��<8�c�N#ya�u��Ƃ�<�.A�S_�-�L�����+�_Pփ��/���x��/�)NSȲEzHeAx�%�_�G�i����{y١Of�����x������<S�.��g�UP�ҳ�Z�}ED�}J��ߏ d���\��'�0I�saC�i�R�X'��[�%�3��a���|j�Xb4�h�����GX6�Q�sZ�u����G\c	_x�������Q/�	~�:f��HG�������� �0�~�����n�0lDF��O�ztN�����ש�L� ���s�Pч jכ�6##G62ȗ��^��!|+AF���0k�=�ܥ��70r?�VU�.�g�C��7[�����>�p
��c����ܬ��X0�U��-��L[�ͷ�� �[�΄�^Lv���0�3Si�����k�s�a�b��	�`������ڗ�$F1ZԈ�~X�
�}GJ���^ <���v-ǁ���p��J�{2�ܭ:������z�,�>7 �"ܥ΃]xXX������+��T�������z��V߃��9iSw#�a�v��~(}}��ԋ�8��Œҽ$޵ڼ�`�?�k�=�,�-�1�(z4*j]�i'�
��l�ҞE��Qc7�C:E���9��wH�ϒ�f?C_�c6���ݽt��Z�d�0#'���IEҩ��cSB�e)�~_W+�B�o� T����fq�}�?��;���������T��
|Z����V�;�<���WCR. �/�J��wzB�~v�G�{�A�M�S!��9���6Ԉ 5-Q؁�8�g;>z���r�:u��ޅC�k��l�/ .������6���Kޱ)��� K<k J�30d�ڙ����:��-L�AC_���b�Δ7�����ќ�g��Ѓ�A�37�;���x����Y�/���#Iu�澒6�m� �婓�n��{k�aG$5�VG6�S��AL&����=�}ʐgf}����_D2��U�s��t��ڱ �|������;�)�w���Qy��R�^�f�*o�S��p�&��!���%98K�yid�����0���}�9��lPv���/-k_3&Dy�,m��y�����.����J��<x �ۡ8E0<�8���W�M��DJ�x5C�����YR���#����?���~���I�����τ�ҙە[�^��;�g-�f%S�W��� /&a��EM��b0Gґ��TG���aC	������zikm�2u��&2sq�Zs7���1�S��������oϴg��<kE�v5�P��~�UYGZ%0�I0�3�t�ŵ+NA�)�<oH��3��}ߑ2�胰�*�2��4��j,�C��n�p�^������E��wS�,����_�^t��H�J�e�z��ժ�HJǗER��H*7q�OF���Żx�&�²�{*�	�w���������_zQC�\�w�N�.\,�U!���z-�����������r:m>�W?�m�E�{Z�6#���u"� *�g�����rgqc�����1Rmeb��;+, �rϭ���Xg�DTʇ��^�N�����x�� ���{��6Ӈv�AFdW�ҫ�ǉ����Є��Θx	�G�FN�����yK�q� ��-�s���3�#s���`B�2���BRU�4v��.�|b"��ct��:���[�_���ft&����g�ynQmCH۪�NJsC5��e���=�9��~~B�]JD�p3��)΢�F�b�ϴ�����Ĉ���"�m�oz����m��FKq�SjEn߻\�X`Ķ��.!�g!�>.�I��T[��M�����anZ�J�	%R�\$���?H64v͹^�C2[;����O'��6iۧg����qJ�Vw��Vu9�ė¿T�	�pߗkD$�&�
�ں�%�,�y
@ֵ���`��}����2(���J}�5�\rB�ϓZ�7�w����G~?O =���[Go�ٸeΖ��/���q��Ԫ������X����W
���,� �|�T�5,�$b��� ��m4��'�B�6��|kp>�
��9

s�O�-;*����7��DWī�<Q8N�,������y�m$�����16�F�j.^���AB[���d�?0X��j��ܶ?�%K�هIw�vՊ2|2W�9};��W�Uh�����5���c�b9T�|�/�':�ً5��Y>S�;�h@�K3����P�-9khz�e�P�&ت�|�l�5ujke����k,`SL\�>������=(rq�j�,�y�z�:�y���!��5ͼ�]�|�I�T��hY���e��q�5�m\>���2�$���!L�.o�A�Q��[v�w�E�`S+�@�q6���?�S�m1��5�<n�uu�F YS�n.`�+��3b��:`^��B������_��w�\o��P]���6Jh�U�`��D��������i��l�/&�Q��'�sY��I���nD��z��?AG`���6���Z�7��,%.��ETk,N<x%i�wd�}K�R���2�6g���d��q07䶶#�TE[��W�$��\�=[�1S�(��	�0ك�%S*�,��%?�T�~��dF�Iޓ�#N�"wJŨov�
T��p���?.�`�boY���F~H�]�\ ]lp��);H����P�X�d-���xj�^�a�p��Y�FO;R��s��+�P���H?R�^h^BٺI%}��q���I���5�%�4����:'v��U��{�J�!���N���j�sr�O���[#:�u�9��x�##��xΆ#��R6p0b��&��o ��7��sQ���T~B�!۾��߳232I#�	�݅��(^�R�`�͝t�%�Д��:�M�c�`u�ĆuQЧNL��"q��ϛ[0<�2.MJ�Yn���D��MF�lv�&�AM ౝ�G�z*]1����d6�nQ���e�	��,�0�nP﨓���qW�w�_v��q��pox	2�-z�`�Z���K��Iw�^�x�z ��>��h��o�B �2OYµ�Aa]�� ���^�� (�r���h=��7�7^�s�A�������D��!��hnq��A��2�w�ȹ7�Z⒆J���^���I'"r�=��W52�.��L�ޣ�Iw7�eP�cj�ֺ��Ꟑ��ed���Ǽ*8�?�5�95�MS��P�-^{j��e�(9Ovw*F�(�d@���+�j� L��l���NbÏ�����Y9Yr�[�&�CQ�~��W�Z�%�*�>����8�˥�_�m��Y:�x��X��lX�����͉a�Vd�)���=��;�]hD����3C��6N��mE���cݚ����\=�ڣY~ɠ�η�*K\�[�(l3��y��7+��?m��5k�s"U�s��|����l~��c��shOx������O<pތ=��,���[�-=��}kb�@p��8�XQ,xC=%�h�"u鿮��L �CǪ������Z��rN���B��	����2kC����n�<���\0	1$�S����8�	���_�ZM�:`ba�<S����h��V��I�[�X�Ii#d"�@�[�hq�c)�_`�;�PLQ�4eT�b����C������F�s�%M�?��Aۯs5V��@��+�\���y�_N%w�c�y�#ɝ+Q����v��%���C\m�7� ��F��TgP�]���Ѐ��!3�&��\����%���6�n�{����A�X��|c�3��p�_�*��N�r�T�Ó�s�ʝ��"de�5���hsr7��qW�B����
�䜴��w�%�5eC�,�[��7��kr9.�%�!$k�G,���2L���F�-T���Gǯ-��%p�~E���bG�2>��ׁ����!K����ی���R�#�$>����
s��aU���:\��3;�p�+�M�������PI�\���A�`"�]���V�xP��H:{�.�@�9��+��,6՞��>��T�p�5�����u�5�*�N9e�s�}�nؤB�EJ��35,��}�Љ9-}�Ց�m�`D`�6�ա>\��%�O�Kٚ^7Rx�/���Ų���+	�1~Ձ�E�&�ge!P��*%�l��i��;�:dV8���Y�©�͸�9edΔ�k�Xxz�m�H��P�>���{@6ڪ���� �C�>fr��ȿ�5u�w�31㣪���ޯ~�l5
���T��0�~�}*�=����28U��(���u}=�]�$0B'�������eQ���҇�>m�c�.X9�)(��=��G;����i?���86SY���: 2�U!E���J��]ʊ��G�<HS5�6"8�׾J��� �K`ia���,_�"�˒�	LS�Le�J��@���C�:��ɐwxN(���j������������d��6��5�*/tk$����[�U�2���D'�e�Sd�drN  �j���3��ƭ��ZǟYU�[V���dT���Ŗ���zI��H��I��P���Go�P����E5K{�z �o#�����M���)�y����z��h#4��#�V���U1�Q/��()����w4+!Q���N���$H��%��-,���:�)�(��-gM(0��~�G���C���h�&7�]M%�ο�����M��iB�|3O�k�Β��nX�^�gp��l����Tx�UY)�5&*]���)z�b/3��5� \����*-�W-�{UV6@A
`���j�/Z#�d?̀��"r��97�� F�P�������XN��]8��E��{�>�b�U��Ҟ��������iP�X�����ϋ�v�)��gB�cɲ�c[X�@���m<r%8�d�^�,�G�p+���+x�R�L�9��Y\}�)�n���6�(b|�E�p��FӨ�a��F�L�8r�τYJc�iրԆS�:���̛5�-/��;���uƷ��\��,W�%�nmD�g�D�<g喆@_p�L}ZTIvKF�H�%ls	4�?򥗂�+z�nAY��烑�A-j��� 9�&`+�� iQ�Ȁ��XH��(~���p�!	���̓�pq"�ߌO2^���!�p���H����� �Z*��c��`����ٿ�P�A.�5�rq�a!.�Y�����m[:J���s ^���WH�g�Z�}ŉ�uqǒ�KH���4�@��Ӌ��j� +K�g��Q_�t�{�AK������X�����S��Vk0�t����;<��!}QNS�eë?u�!w�Kr�X�Qo���n�@wJwh���`,n����-ݯ��͘�,���²�{�X�MγS��
����$ݤS#����������Ջ��L
�򰘑���ޞ��@v��l��k���R��%���mq��!��n1��խ!N�ځ���r���ͻ���
�9đ�Gi�bT���s�,̚ld&��T����F-���x�K����)��!����뙓�Ή.ݐ������VC�ÀB���nz������	�v�)./�k��*�I4<Br����;�9E�_j�M�NZe��y�&q�	QJ�B�A��RǲN¤�v���HvV0y�p�	�.n+��t�|�����6vI�F3�G������^_�3��0u�<A�H��-{����l��F1�(r�c�"���|�p��?�Px��/� $1$Vv��'�_6P/k&��Sq�i��]�M~�rɅ�����k*|��R=�X�i�HfA\�>%=}�G����4m"��̑��%��|s*����n����wfU�x����G$(�a��*
�0'��*�e��H��za���G ����dM��D���㸭'y��t����3�ZR��g�����tr��1��]�	Q0�yڮOu\�%	 ��f��<��ERr>p���q�B�N��>�{�XU`Y�N���e�Iķ��Ӏ����i�K����w@��t$LN;h,z���¢����,`��)��3#-�90A ���y�1�Us��1O.�R�YԎ��\�A�����^�c��.i�T	�v�Iʰѻs , �6��=� u�Zg'���ŗ����(�q��*�f����`GPD�O��B���QL
��^�@c��5!���T�Q�I�]�2B���j+E��}
ZSHAy���Pk��Ҭ�w�ji�g|��Y����6�Ҡ�8y�w^U]�ۚ�y�Nモ}��ҦyT��T5�@�`k"<"Fy�fW���P�#|>n�X�d)�"JF��4D������ *���ʳ�t�J��G�D��\�
�v:dw�Q��⭱��w�8A��A���|5ғOŎ����;F�� ��������|�;��]��ԙ#�<�،Խ_���|.��g僲��<���5�z�bI��*X��=XF���h�C�D�"8:�S��V1셷�db�ðt��6��]��� \��B�P�WKX�{��,���a��]��:�`��:�	�Ö<3蠜X��4�u,�s��?�|������r�?r����d-O�=��+&J�}�O��$V�
*�M�'c)q }+���rE
��Gӓ'�^�L��(���3�,��md�5%ÿ��wCdl;�5�����8'����

�ŨӤ�J���B�u���$F��|��9����N�<E����){�;���]���)p�/+���L*���~�vA7a�b��.{��3T��� S^:�0�X/w�="T��loV����R�4��" �(��_8Y!=_��ȸA=�zV��D�E�DѠ��B�Zw���)tT4`홌L&X~����Oj��p]�����V'IM��u�[���@������죹��MdE:�P�<�*.@����o�����ʏ�;��(���7uO��"�\���|�9�V�+:�!e2'4�ݵ��_�C�	������5 ���M�D����I����!�M<���D��Q���|�]ԲB��4���7t<����q}��n�ӆ�1ul�}�ܫ�[�3lu���s�E'���b�XY��|����� ���}�%�%�����ϑ��_^? I�B�^�Ҡ��ſ����Z�bt���� ���$I v������nhL�/����_�tNYČr4�*�x�����;T�tQ�,պ��*f��ag�M媁�U�8�(c�K���1��mY�Nf�Gu�{��ר"�-�D�)���00��0��rS�a�W���33��l�K��'3��^n�`�%�T��?���|�p�y���~C������"�4���P�9r]jY���>����~��P1:x������� q֬�r5gYU�2L�����Lw}��W�	���b�n�dN�v�&7� �-���
/�y2�*mj:BB��%��N0-�.-�V,*tIr3�,���U��(!/ ��?������]��6u�����^�_��-��Uo��`�n]�e�أ�x�-~�#�§@P������b����op���>J_�?�%؏YL.�o�b*[��<v^�P���.S"�r��kI�S�O度k�(d�|U�(�I�l��ӊ��b3����JӏR�vA�VG"����O%h7( �1�}��N-�m4~��s�&yd/�GyWV�~P<���)��f�G��W�f6�j㿀%��j�^�Ť��2xI�cGZ�I9|��v�;=Y��h� Y�X�a�2�>,o��K���ZBw%&������'mŪ4(���uH��w�z����ަ-q@ZK��DPP�0j�qί(@<#�C2W�h}�j��p�m��4�]��x:�v&�`0Z|����>�'��~���|�+1���3��,!
�*95gkl[^�[1����b3uD"����.�W��Q�Y�����E{z�mX |zl���hE�" �L�I�X�o-N��%'�)%�B��@���Y��<�N{�qr�wd>��Som��`}Wq��O`�i��Af-�V�7{���\�P�����g7o�˴�z���lB��0��d���^����K���tR��k�>�q�l����x'O	�E 	<8N�o����l�B��s��F
ar����B$ P;�(Q��s��-'a�$��8��01��t�����T���v����}���O���� XE-�E-�F!�Q��a���^^s�<q��k�9�K7�VE����)|Q�����b�9Ι�?������
���'8�U��U�;!W��\븇H�e"��x�u,8�	� Z�Cؑ�ʤ�$!l,@oioa��^B�+� ��\=�˸�2�$7lqjvUp�QyS�l
1�c�Tv�b��@�!B�
m$�z��-m[c�H��Zd��0@bZ̶3:��8�����X�Ϳ��#<W��/�=��y�BQ�Nz38-#�3�����$�i�(%���&�M�=�Q# ���^)������)���\��J����W!�>v ��.��4� �'�أ�ѫ��`�C�������iA(s���.o}����^��7���O�v����A��!M�\���v{sV~^a>ԇ���N�Ҍ)��A�����ΒL+;k���/ܢԃ���>�j*ۨ�eW���Ej/.�����[�A�5/�M]����\VxTՐ�&c�DC�c;��f��	�d��!��i^mh������99�i)~6bD����Z#�v�A����X���ja}��U���as;�0Ke�$���~��F��q���C��1z�YR�;�v�K����te���Q�FFj���\R���'4�sZzdni5����|!�p�2w`S��y��(T, �03P��|�r��"�m���컰n�6��|ټ�,��9�NM�Fzi�>8��C�>��Ţ}�4f�BD��<�czף�=���R_��P���v�y^�ql��o�z����������:����Cr]-n�{���u���-\��֞8��R�^(^J
)<m�%iR������@����m�c�#�Xj�T��I[���3yq�W������%`U��`��{;�������0�a9+2>!�&?�4٪'��A�q(S�nP;��YyQ�G�HۙG�2�(,��dӠ�@�wDH�2a��E#RoE'u���v�o�Ju� U:/}�7���<N!������T!�*z�tW*#�H5��>�����Sb�/�P�����(�6�]�d=��s��8�jbꟚ/�!p���$4/�����D\���ۍF&n��}Oe����WXx��������"S�ㆶ�F�d�4����T3��Ez�Lpޣ3c�ۄ��������K�i�[<��=u?*�N����5�4��ВΊ�=�8��J�H�`��G=�#�����	0�l�M�W�,L��r�?:qu�P��6�$��
MX�cH!k�ߨ��0JX�� ��
^5�{U@vצZ�q4�L���]>��Un�YŅCp(0iW ���~���p��7��:6k� /�z�;�	�@/�p���4�k�B��-��N�S�s��ܲ��GuRGF�{��'o@��E(���R�{+
��F͡�`Z%� t�%
9���Nk��5��?�����)(���W"�H�--�?%g{M�tֺL��!|���$QN�8�����桸��z+G��:�%�Z"rխ��"����ڲi�N�m��5\�:Ud�Nt�/���vX��Y��I�@'�?��Jע[�~�Õ�{.��ғ�Z����;_���ni��JRݥF��y�po�-�k2�֭��3����2e+)�'t��tT��U��\VBqt�	�^F�۞m�U�������1���J�hzI�$�JFMa"B��s8`���oy�X1X<��q"���!$ߒףG�)7�4��c�CEm����������M��>��o��w��\C}��#QP��;��f�!��`g	'��%�vX�}���.�zfB1��J�*[tMa1�1�)�C~��o4�@]��>s=9�%2`�Is�Cl�]�[ m�9e�-�̆�Y�MU."���L�Ѯ��|G"���@�&��������D�����4��8(��(�5#V��-+����/Q��!��r��f/�|�%m�Ê@�o�/ 61	�":$��򮛼zW�>������rJ1��0Pܿ��1�,6�n�Qt����?!�iͳ$08h�~1����s@�<Y7��O��R�~T� �o�䠉[��~{^��T����?*��N��JP�ƾפ*Ms�Ek���-����,�cז�Z�+�A��[,y�h���r����a��.+/�6�2�A@&�NOK�����/�9~������C�P��4��Y������d�Zl�QH<�ɖJ�Dۻ�}y��%�})|$�F��� ��d����4k����FvqP�<�!�VZR�D33��գSX���dJX�S��U�x��lGޛ냩_Q�p���ݴ�P�M#k�6TBg,͘{�	��ւ��M�����T.��{���1�ΑثY��a�xK}�_Q��gQl�X�Y��[�h�q�-w�:w�(e�=�w�l�	F'EγEݘE���N~ѦUõ큥��w��Ofh���[M'zÞ��<��}�}�o�

VP��Cr�`�un�WqX�?����N"ڈ���
�8H,�aD�u�OO�0��0��cY��@�2�"�\��d��D��vA|�D�?Zǫ��Xz�d�N���������W���:�]�>�����cM1M�@yy�����*�m �:ͪ�sCe�
�0��[�� � 2��OU�h߇9�VH��Ѻ�����r<��-�Mle�r�r �y[���N
a��	�v��G�aDdǽ��|1��O�=���+�cdt�|y��z�#��E�Ԩў��@\�����5/��ʏ��'��*��NH�T���b&W�s�([��÷�1�xA��(;NM��+�7F����(B�l��!AF���G�g���id�۠m��"K� :�Q��N�f�����径�9Sn�D8�����]H�Zv߻�����7�'�l�t����Bs��2�({�����V�K���c�]im��V�l�4�r�p�ýQp��X����|��[a&%��u�sQ��fc���Q49�������Z*Zu2b{1�j��`�|lab|�*��Q�����ӯ*Yx��Da������eH�i2�r���3`�ߊ/޺O9����d�f`�|J�J>��|�#�y~�%��:E}��e]��@�����*��\�&�_%�L[b�'�"�\�Zd��T!9]�o���>��D�� [����_G��3Ƀdr�X�f9��n�mk���`�7e��6�ʆӜ��L0�t ���
a7��A��D6'�ܪYA,P5���!��4���a����'7��f��� h�Bc�[�\�a��P:\�J`U:`]D��O�m�XN��{�`���z)��Z�y�*U�AJkaa�$���� p��o�|*Ź�s�<�>8��B��9���� ��Q�P�b{3�	�>�y�D�Ā���߭`�2^YFi���~
������d|�!�_0��������dG�=�����7���_�B���&Z`������k��Q��R��AMU#�.iq��B��\�J��|�6EgA���r����Ո��ۏ����M��^l��^Pdb�Z���+.Fn�?�Z���Du�`B;��姎�Γ�E1��Is�8j�a/��Vq͕"C���ڤe���<��!#Of�v�)��XF�/,+�8UbH��8$=��&P��
��{[�'׾i �ʡ��	u\8��H͞�8J��FQ�Z��������6?���>�/��Gnۧ�F���+��L ���;��i2KS�x��9��]�ܗ}�U�����o�4X��T��oI���$| oHnO�A��ЉUȄS�*:�w�P���Ѵ�GShq�l�.��L���ae����&t2��xT#���<��d���>W+����f�95p�
:����mu�nBxCȑ��8is�)%�GXB��/~��Z<�������qt[��|4a�}��t�W���#���H|!7Cf���9��,u·?ዒ�CwU���af
1NL��&���n�?���Ǩ��q_�A�O��F�=����Ux Ѷ�r&z	3�Z\y��ߋ�,ye���M�q��E�Rr��;A
��)�P%2�y��I'kg��M�VߏÂVs��v!��op��HPԔ�Y�"��ӿ^&�Y�C�U<:f�w�_/J�I�T漾�i_�$V�֥�/3�T���}�����}��8XQcst@���\]j�/Ӽ���5��S�O��F�G����3��[V����^�x���P���d�����iY���_�|	�G�g�}Z���?��8U� �LJ�xK��)
���J�%TBa���x�k�Hw��{�ص��?�i ��s�3#�y+����gZ%�d�7K�߼e���y&)4�▕������{�c��⼹���ڍ�@v�:V�A��?�'D�:��x@��ڈ^��-|���9eH��*%���}<B��g$���H>�7$O��L�d���~5�\�gs[ٗ@I?s�rf��`�E��&'�}�"IX�Q�6�ܢnO�K���?����s��To&�����eXS�N�\�`t	��w�,/�[�}{u|e>Zԁ�--.�); ��t>�q�m��k����`e�����$N�=k�\a����,�S�x��|!����`�_��;�H�>�qE��F�Ҳ�](�����S  �x�!�9�Y��ǈZ���m(	6JM���N������ވ����쌽�oP"��Yp�y�s��h�s�j6�V̻э��bԃR[�����l������!���J���|��t���2��oKggvK��L�����J~��G7\�t۸�M��e���/��.���\��Z�m�;�
=`�)�z�AvDUdpx���6�πe��|�u�H�{m�e �E'�N.K���<�T�K�`|�����i���Y9&]ڟ������0�5+aE���M7��2�x��aO��a#zt���>���CFKT��8Pi�&����KY����S����߳�
_eW,�N	/^e��Aἡ�����z�(�5 ;Rmx�."�	��J���_hN�u��THJ��r���ރ��~�l�d,�����<C�
�Ȋf�s���8D)b8�>D�����a�x�kV˶������T�ע`�d�:x�4��I��A�l3�=X��[�'�n�M�� Q\`���q�)�����>�;�KUsLWё�w�ąT�Ws��͞��� <����mcd�_��זz����Zl��#��c��'�P���&�{7�p{�$�1�k��~$����:��*$[�X���G=Dk��D]����5�����ZGZ/�q�Y,��q��Z4�:�I�_"�JS��?��.�f�5��}��=m5b�J�`u#�@�R��YRBg�����@�c�e?NP#�e�W$x�s��M�ɨ��J��5�S	ꖎ|��Rb|;��^�������t���H���d�v�����R�3�	�����Q5T֖�`��"S�Y��*\�ȫ���c�]�Xr��M������l���I�(�Ş�1��	��:��ǜ�)�G�Y���'O�J���#>��6gː%�nVU��<S������6K<≾�Hv�&�=�.}[���(+S�����A��	�9����%�]|���]���WM�tO�ȝ�!#�LW~�a�./���3��QȘ~��e]-� :bcUy�=��R����*]�߳�����O!��)\�Rp��]�Q�R٩��IԴ�h|@HR��N�CF�;�荽?��e�,R�=��U�7�l�K�L��˻x0����|��ă�J�9q�dF��彺��^�~*2��L�{V����'�����m��S#0l���|x����`.���L����+�slI7���(qN�5�i�;�N��% �9�{M�����_^W�*��p��:��^_fX"�t<�
#~G�v+�#30�.ƿ����Q�^��EV`?Oe��l6!A�@�2�6�(���G��k�4E�p��e)\e�h6BSʰ�`�u��Z�y	��UmZ�\����rRp��q�"O����s�!�h���`g��'0rq��3a����n*��J:|.<���{3+�G�Ja ��ns=GMz����s�;W=���7X�.�#��N�N�dM	#�܉%�Y�>f!�!�֞h[�E��`C�m��z��UH�=P�V�]����Oy�n��]	z�ͬ4Fd(Q�U���}�P*�#��� �tR��g�D������=��Iل��ώ�~4���SRZg�Zbn~p>`Hbвgn}��$ͪT�dbFH�p��#�h�ϱ=0�P�n��<�>���u!��o1{�=����L[)dx�h���z����9�A�]x u|]���m�@oc*)�e|#~8����"Dt��|iź��1�:�#;"���G��Ik���UN�FsA�-�X
#Գ�bCy��'r��!�����5�o2^��\��%�hr@D��S�b�
��T��3N�}�*.8��Z��4��-�&Z��;�����&9y�(⣌,Ҕ"�}�����ט�i*�]�0 ��.�s���t���NH| i/�a�W��T�K!&�_&��1++�{��A�P�Qo0�U������kǛ����L�f�̓Cb���t���Z�CÖ�i_V��/ֶ����N��5<�J���=n�Q0Y��f ��AL��|����z���=����$;��%X�/��z��a��z�i<��l��:i�����#/f�*]^��V�1۾�pu4t��
}J���db��v�
|<��;J'�A%m�O:p��CG��`���\�����|���Md�_1_/u0_�{d��}���ː!�L!)Ͳ�P�
~���zn��2��3V����N}�]��$靀y���q��s�H��&G�#�R�`*}�2[�҅�:�h)J�&��D� �\�oc��~dVLR&������.���=ɳ9G<:|-a{]���R:->���"{޿�7�+䯊�~#n��;_t�D���d}�D6d�cW̊MJfQ4m{s_^���j�K��g�f l�S�C�.������wpuR̅!��q��oū,�ODj�j:+iT(Vшtt>���$+0غ5wH� (�.�ꢏ��fUK3lƩ���XI[SS��n�Nc�BVY�0�{4<t(����L�{��_�P��:��%3�ݸ¬&�g�ӚR��N9�|K�Tq?W@�sf�s��ʪ��}�ӽ[Ĥ若�vw��zީG�3Ge밀��v�F�lt��嘪���� Vӓ~Wa��]2畈��Y*"�m`>^E����>h��bT<R�p[B�s�EQRC��Qy+3�R0���W3Wߙ�O���2LH���b�k�K��!��cΝ�b�Tō�Ӌ���<Ԣ���x�֌n_�Ǡ �8���"�l��l^@����8�na�\�iQ?j���C [!5��o�SK4�h�T�z}ߓ�ϝ�B��a��0�E�b�HG�uq� ���p[�N-����}І��I�F�)
4����b�s���!�B��}��X�^&?�2k*КWU��rd�@��a	�E� _�n�R��/�:=r+m� �?��L�`_�P�$p�s��PYi��#�j9�d����a���Z; `�(��A��L�Q����D�$�)H��<��Uz�-�0M��h��e<�J�<��m��N#���oW*d\��?bu��t���2�x����~̎P�~����l�U!�pˇn�Y�D��^.�M*h������W7k�R�oKr�C}A:܉Fo��c�ʹ@��cC��tp<��UV���#3�ݿ K���~U^f��b��y���r���=�K�JR��/$��^M|��+�n������d���l%�^\��l{��_���%gt�ꀏ �]r�iu5��МR����N�I���T��-�U�ҧ�Qq:
���s���΢�:��Jw�[}�C)/�h�I�Sw�c1Ca���O:K#��T7���|f��o�u��KMCE �D�&e�
4$J/�B��b%�ֲ���Z����}X+��r�Ѕ�VImȺ���T5+�6@ѭ�e��L��vj�o�k�oB.�T/9���YT�i�;G�/�R�a�A0�M7�0����Du���?�sy�Z�n p������c�Vc@(u�r݆�AǪ�^��T���i� �X����r�S�(9>3�<˺�N�-�l"�[5���ǉ#�Q��ʞ;�LD��dd��ɖ�D|z��*D�>[�?�E�<%)@�r	�� �+�΅G}Q�DVC;�t��=^8��,A@��֠9�iƤ�fp���^���!�6>m>��N�Mu��Np���`e:R��Hh��wU���{`�����3�~7�p }ܫ��x�j��(���x�1{�tU��{���5걐�����Q�A筮�=�fpG�;D�l�c�I�7�CV��N!�p�>�r��[�U��O,;��ihvQ�)���f�&x���úN����à��no.�}v�osHt+~��L�2���Ҿ.o��3�u�m$pdn	�C��2J{� �Ӣ>�Of0('�!6�I�
��DФ!]vD���{UBv�(cb�P���3�*��I��[�@�bZ�9�d�}*X�`�3Qť�kN�:�G�Ϣ�bw�+&n�W΢���3[��߄��%Z��#H�^ޡ/����Y�1`���%����j��p���\��bD��3���vw������0��	�u�� t�
���X�9����7�j��WP3; 	7��4����Vi&��>3�
#��UM��{���Q�m�Vd�sp>��N�~����uI	�{��[�܎i�ⴜ��)l��c�B�)��C�f_�u5�W#�NK�H�a�D���ު�+��żߡ����`�먋ߛ&��.�Y�fM��G��zG����P�;͞o���c� �!w�I+��&�lŀ�� �3|����(���l���
\�.�����#r�%2�h!�i��w�$p�
 O:;�f�d$aKg���d����C�Pd3d�+�C^�i�5}���;��>7jL���p�;��_e�s��?�K	w�U��[�A��w?���m��P��Ƿ�Ϡ��R��ᖎ=��R�~X�K%��t�S�N�C�� ����	��6�U�;o[+:��ѩ+w�	�QΪ��c%Oru�:��"�lWs�ۄS�Kͤ���D�[����Ts~o����X��gǎ�������'c[D�5J6|D{)����Y����t����w�����A�?ER7��-;��hǮ( d�Uδ6��8N���:G7�B��$�5�69.����Tq�H?�{���0ڭ�K"�z�Q�,}��NC�ĸ@�QF��nƥ!��S�Y��V~��{��������`Wr{-����|`X��JjC�@)�ȵ�\ȠӜY_Ӏ���8�zVn�}�fί�S]$��%se�����!Q`ֱ���ZE8�xُ|ed��j�7G�H��r����8��NUF�Ri�z�Ya�pg]�(��dLM�q����f�8Y��7iXڦ�sǂ�zr�`�'K�N�
�a��Q9L+!+`x�<�q�P%�WeΈ��ݺZ{�-���d��>���V�}�����"+E�m,��(rb�f���ɊB�"x6?ݙ��kdi�]�܂�#��d�����@����Γ/>�	���Ӑ=k���;�w�E��%^i$s�0�82��� �9��,8�?�%[����dC��x���sb4� ��q��	Z����K�IV�q��3qwgFJ�l� ՗䆻,��s�q��Q�c�Pl�� �q
���9<��v�(�J��H�`�����'��T�_���5Y��0��r;d9VBV�B��F΃���ǌ?��?(���VL!.O�m:���[�t9��$�֟�C��0��c��v�M7\+Q����Mb���8�U�"sz��M�W�+�싆M���񴧰Mm�vئ�C�8��0C�+�i�oj�W�p_�@F�h�9l�&�&x����'gϮ�ҎUs{}� �&�ץ�%.���᠇T!��&Q��d��v�mac��Q�/t�Wm�C��'wcDf6�оDF�T~W�͚�:E|��]�!�&\J��,����0(ol��B��� ���D7�[����Hj�왩�鮳3q�6�Z��՝5p��YdIέ8�wϮa�5�u�@j����.���v}��ΰ4�3pnqx��� G���V��L���o&Z�Vݏh����r(�_tp����Jpo;�Iw1쐵�2Ϥ�H�[bp%U���*�}�r�	C	����ԇ=��k ����ROS�G��b��c0	`�oI C�Y�`,���|l�Dw���j~�qF�0b+�Pf���L�m�+K{�f2��C?�a���D�ğ�px�R��v�}^=FƢ����y1���V�M������+p#�l���{�02���<E8���{�hw~����������#�s	 �����\��S�p;:��*����E��Ò�E\���{�^R�]��u��`,��)��C�5v7�.n/�
���T?ZT8Z��V]��<樤h�!�~��ǵ��'�'��Ue�ԁ���(���A�M3d2�	sX�\Vwk0X8��.s,�36�|u�]$�/W��l����[}��'o_��m��XRy���_�Y�66Rxaj!����-/���8g�Ґ��lM\A�Q�_t�|P�(%�A	 獛��Ə@�s�7���#��=G$�T��1{�����%�)��?�e��H'�/&��o^Ȉl�!/�38P�;>��@��z���X�$w)�(��W7"��̛U��X���Ucz���e��"��5�k*��	��AS���3�ze}(z
h��*�)҆�51�?KԀ� 8���v�(g%�,��awG3�iDkK�.SOb]4����2�	+?�զp?�=�ɾ��D*Q)@��]"�{J�J��u�e�c��v:@1n��-�4m�ӷI.ё��pO�`)���ЦaR���?S&U��nZemH�ɛ��B�R����Is�K���"}ۡŶ���h�eqH�,���f[4բ�7�ɽ7*���c�!���b�����
q�3���Z�kˤfM�|O)2"m���]����KKGy��N�G�B�Y���Ju�瀤U�\���1H�-B&�c��ǄN��ϔ\�e�HX�];��>ʔDǰ:��\�m��oڿh�ߦ�%g��٢CN��E��OGL��¬7Md�3�B�O�N�ޒ9r'�AխQ�%��
�%�K��r�����͗�}�|En��Iʂ���,>�W4|�$#%�y���LmF���#�a9%w�%�h�!�J=������s����_���3��]�;0oK�'�P?Ი۷��۝�oº)щm}��|�,��m�T�Tv*��M��{7���E��ۍKI�>���;W��%v5����V
XW�B��E�܀?�]{����4Vr���
�Xt��W�p��j�7Qq���Z��z��6�!�x��۠�U1�z����+l`�dsV���,���̤[i_�����-�<G�� Z���H������[���$ѿw۾�J!��t��W�������mT&���.5;6L���u�p*�j6�鐉�l��:�)���F5�#ܥ���Rߤ��S膱�6��6:)L0���u�����计;T�\āu�B>�a�9��OD+lx�)�k�PO�"�_��ǲ"�y���O�{'�nrU�()��=aGj(-�ܯ_x�{D�iq��iTp P����BՐ���Z0��Enz�S����qU.D��r�=��f��cGP��EŚ����ld��Q���=h��)
������X$�j�nLKw�˅�^Y�D��t/���NpC/e�<o�r�� 8�K��ITa��[J�/��eJ)9�L�;��7Mmug��gϞX�s��C[6*�����յ�����$s�'���Cz�Mn��\	�ϳ�ԉ+�*n;��gD�3p��#��6S-��O
�y(H�;��̻�?g�p�k�и��� �����W�i���,q$K����x2�i�%��mC>�Hܜb���Oٞ�D�����5����T�/
�"!�[�9!�R^�̐;���$��Ìh
�p���SQp4n0��=^�������rx�ɀ��e��l��Q$�m���ދ!Wѧ]U���x` !�� Nmjq��=�ádz�J����1��i�+�s��fR]���k"�&u2*�_�����m�<��DxE��ה�����I�F���,��]�4�R�k�@ш�$ZI1�n�}��$\6!jHhA-<�9�ub�oep��v���v_��C�қxU��Y�	�|]�)
#хr��3���h$��;���-⤥�%�QK�q��΄�S����R�Ƭ:�4���|d�[.����X���#�*Ad�	з�����nh[bkt���![����q򜽄<�`��Gl��y�l+�ᘷ/Õu\�� 9� ���>��L�t&���wz�3u�7/l��B~j����@N�˲S�tJJ{8���V6���č}���H[�"��0.�u�~^0Ƹ�a�+� d�po����zN���7Y1�Ӄ�u���W���R��f���5�>�����H�;�1	Z��a����v�V���6V�����	2�<؄���Հ��>���Saz�]�(�2�3�X��L��H��;F�}�PG���p�16	��u26��q���/I�M��=MB�ty�_^!����K�d�� ���`@�P7��(C��0��z�4M���\�]eۣ*1�¨�����Q�Լ,o��بH���S��i[0w:��=kz8_i�H�Ȅ���G�B�BC�cA���2�Im���9�
��u�O�5����D��2�1^=ue�C4�59VF�qy��e
VP�v;�v孱���{�VD�g�4 ���ɘ�*]@ӥ���A��yn*� o��z�3_�4"�*\�z	�D��;A��_Z�fޑ21&��
ΞG�]��r�A�>t�?�G0B(��
DT�{, n�,w�By��-CSK��Ѣ@��f��𾀺��f�\Ҿw�'���pH�J�'h�^-�����m,� J��J�׎X��(ǟE���S��\��Qғ����b1�if�R����÷J�-�E�΅���7t�4�@�j��EZ�#���q��?��
vE\��	a7]�����G��Y�M6`k@�k�B���!��1dug���xj=�ұ���Y�S���9���6(~|U��U�;�����1o�+K�:��M5�(�wm�Q�e��Y���h����Xq���}�M�u�p��f0�g��x��i7sE��Ͱg��D�c��L1xq`�U�Y�&kva�kA�>�φB^-D�2EHE"�Y���⟈�S/)���8X�ѭA�L�!��R�/��a�0}��D�ۇ&�� ���%/�=SW�&|ky� )��Y�ѓ������#������+#�{��"�Gnݶ;���M!4,�!��p����:��l���ۆd��r�p���xۏ�޶��J_�z��{����b!��/���Â��I�`O2���2�7L[V[�v��2T��\(b7�喕
>I &�������~�$j�X���@����.��,jk�\<^��kE�Y��.�t̄�#{8�9�7��/ӭ�ƥ4UpY��B�������J+'�<Od�}z G@R�����2������FÔ܋�&�d
s��=�#��dJ2,�#��S�ƀ1a'S��N�L�OD��m�Z ������7��,����0K�oc��1�jd�:{?���/��E%���ܛ8���w.�^�T�!:y_ٰ|V���v�[�5��{oݗE�h�@GΪv�h·9"���˟?�s�ն	�fY�/�r�\��xL�ٖRQ� B�*>�A}���W�^N-8jC�_ ѵ��Y�\@��ݾV��ꕪ*�����t�c�n�Ugf
�;����%��t��p&L�3ح\���cU/�/$�`�ɰB�p���:e����B����z�0�+k��0��i���*W��<��a�t�>��=g�߯�><��H�5E>0�`w�B�6�5@z�c �Q�9�L�k�Vh�0��+�t���S��y�޸����$�
�������tc
Y;a*Jf�їQ�h�T�&�L��]��F&���JJ�Z!g$�X(b�*�4d	�r���� �h�Sl)�1?��<����\gIx`+�\��٠�)�#���c[�Ҡ�'>㹈J�7m$��Ǖ�r݇Akbsb!���:S�ޚ�
֭�^-,)�M4�>��˔�`f�o�Hm�ꎏ�C_�v�v����1^�%�S;�ڗ������ݙ��&�"�L�gl��t㰀�i��X)T$�V�wVG
��)��H���t>������VI/�j�K}�t]�b���jh)��d���թSCK��NF��¢�lAku
�	�qӷ��A�?X0_Ɓ>�ٖ�����߫��^�]�meD�
/���4,\�lt���kx9W7��^6I �P���p��OR �4�_]�A{� l��V�~�q�����@K�����=��l-g�6̝ �51=��
(:xjѸ�nD�Ҿ�!�D�)o�*���:w5
%����:d�\G7ۙ�SP�K�g$:��s*���^��K��5�h7�j�CĻzl�R9��q���"�1��Zw~Q�7�DU+�3���qt��[�ڈV#T�eC�e�b<�QZϢ4������,�8\5��_NF�w�^W���'v/=υ�M��.����F�a]8ٹ��W!� 65h�[)\ǏKF�`��d�b��1{�05�Ə��3�9�~�Ӣ���.=B<����y��ѐ���spR�M�\����r�:��%oW�{��ͬX�4��c���ǧ@c�
����e�����E=i�m�|��A�A��%�:{o�����`S���)=��4��8j����y�Rֻ9�1}A�Z��!�U�|'�GZ�Y�g��u�8ÍC��uz��f�!���{�U�&�'�ԫFN�2O����(���r�!�?����k����k�ᯫ�d"��
&W�R(���ښ��J��#ՋHR[Y}��B<[�b5�X�o���ԉ�}�B.o-)�܂��B�ME����x�8W�����8������x#\����1�{�p@���q�,K5E�<��T�e�ѫ$*�xF �0=��t��+��.��ȏ�F�V��ʊ��bpI|����M�%�	c&K���hn	>!�*�d�BވN�â�l/�v��<�p�x��Ép N��-c�a�� �Z�:B���>L�����lf���ëau0��g=
<!z���Z��	�b	lB�J^���q��H,�	���>�����K��c�_8��1 ��z.����2ͅ��,���'ȗos�e�g5�,�����߅�&�3:|*Ώ~�t�\̣�KB�!�f�:����i��_���ڇΕ�,i"�+T�b$�K���pt?�XU9@>��<�MH2~��1	^Ն�E�T��KmV��g[���6)Н.e��g���(z%L��D=�@��^�oỳ��w�c̲a]uuT�\�������f��e���E��N�a���!Ii��U��P���(,�e�Έ�ڃeA]��p!�Om����`w���dIޮɽ���:�Q�2g��.*�>��V������	�2CҀ�-c� [�{��[d:ez5��Ow׵�S%p�lۮԊ�Im���:���z�}�턩]5\N#A�Hⷝ���G�^CBs/΍��cP{v�%�8�4�bL��`�yG-A"�� K(gl$�0Y{N��\�~zr��rKe?�s*��;�a�f ���	%�vS(���&$Չ���;��6/I�?8�צM��b���)�"�X��C�V�?���P���π,X�_?�3���4��C�%6V2��U���-�/�\N�g��l(�R���ѹȳ�%�\��,��#�sx��ʗ�6��_m(d����3�/!��}"�E�k�*��{m����g-�.�������*k�?"sӞ���t6���p�Lk48���<�5��a�%��r�${�w+)�b�G���tG� � �v΄qR�{!X�˟U�H��@ ���~1e@�F��a���SC���uI�2z��Y�+��m2ktϭ�>� �����U �|�2��&���;���b���U$�<�ӵE�Yhb]����g��uh��+� G�M��Om�S]	�>�A2@���q��R4'jB+�p�x��� ����xm���t��F�v�C�R�J'{��]���ev��Λ��iV�.J��{m��sŷ��.��΁#�Q ���͎ɏYl۝m8��H�jҩ�9w�@[l1�$����*"�����.�;��<���Ƨ7ٷ�7��N���}�;}I�G���%yA_^z?�9��/��_˔5�(B��
�%l���b��.1�g(�.��߬���h�s�%m�� ��\U�7ԁ���c�R��_1��ʘ�7n;�����Z1[���G	�{�v�?�1��렺�	1��������;,�?=3��)%oK7�O6	s�՛�{C8˫��c��1K�<.��Zݷ-���P8��Ss%��ﱮ����a--tCxT�����]5bi��K�qd���)	�^A��tƇ��	��z�3Ґ|�
�������უL8�aU��LW��=�z�
�k�����>X��iJ0�Dws��g{8�T�Vk$�ߐV4�e���I�PB�_��̺������NN��K�c ��V�����&us{�����ɱ?���	[Y���F�fZ��+=��{��^ h���-(��͍k�Y�-,�J���=uy�oE���=����ּl�J���.�@��k���#���b�EN2��������&}��k��<l�E�e�i.K���s�N>��jy�	Ns;/�_�$,����yj����9r�
`�

�2���h�ʧ6u0�?n�0I"e�F��U+,����=A#ɔ���X:�܁�M+6�Y����h �~�`���Uu��ܫ�4$����]o��aH�i�8ٮh�,�Hbg�"+��"�_0ȼ<�o�.�j�aG����h��y�9ț�5�]��6�-���K�Ӓ?t�C�W�!{��+A![�A�,=m��d�|��b�-nc�F3���K�]��U�k��UegQ�	ʊ�i�{�����]E�bE�����kǡ��vfgΧ� 9���z_^>ˋ��ح4�m"ɖ�Uf�Z�~�DNV�L����y���L�5$}6g�w�a�_W�&k�
�%��d�T���T%u&,���%�lq� �9�պ�p���})M p2W�/;R@lel�MHiQ�����-1xk?�7��G-?���/u��	v�)��R`�����6|Ct��1c����|�4�WA?�;/,�<^���дJq7��^�1�|.�D�MA�*�8������-cP!1������;����
4��|�&u�b�@���a�|:�ρ�(a6��Ώy#)�vo{I��I����F��;e+��A�g����S��}I����k����������)�t��E�7����-��q��P�����D�Sa)"4E��U���Yr�����'jmⴙu���\H�w>R�w.�g���0
6���쁖NM�e����˚�k���I��M*�k�q����B�{�h��WW�����w�G�)��g252>���x��}�5|P�~�m<`����&�JS�ĕ�<��yק ��?X#���	P�5yX���;��U� �ơ�4�W���$���+�G��S��:y���n��7��kV�S+�~O�+�٬��w6Zo+�Yj�!�#R����/��O�G_s�cZ?8�w�����	���ZyZNy*E�ʶ���.��8��<���1�WQ2��+t�7�~�����L	œ�V�7Q#/0ҍ\�<&���ӕ4�և�3���W�����Ԏ��۔�&5��p�f-���u} C�/���� S�G�F܋��PT�9��T�F�iLh�����.ృ�6���3�?�42=Yգ@F���n��k��iBK���h;1�նaj�hϬl�gn�5����}�:�cE��0�է��7��pP����D5�V�� ��3�AOhj�bBW��@R�qU@m�~N	
�ݪ��3�i��e�DBX�I�Mٹ�CRɞ�=hjq��}�3��w�R��|[f��yl��>~A�4]fkT���J ��"��*��H�X��Զ0�Q"p��Qm�;v�e&߭A ��l���;V�Ym���hzb����X�{�h�k��'j����v��i�w���&-|�?ˢ�G���	j������'�Z{l����M�x�� +Xl� #��
.�c����\Hg�d�sW��i���Z�.�Lp��u�Rx���[w�����>��ͥ���k?;�w�[쾶�HS�kS��`Іy~�ܔ$D�
���3��.�G��I�����Qw�UX}fA��6�S�3J�t]*��Ub��}��d�rX�.w-���,F�#$W��,n�K����3Ű�IK�Py��z(UR��X�y�fM}V�9�'�G��ٓ��C�,%ڄ���s���T����>F�E��ݴC~�Rtr�i��zw�Ё���J�Wj#�ܭ�6�3m����Z��
���������Z-��(�2�a�xq[#���pN� t���B ,	L��s��9?ly���5e����TF8Z�E���!l�����Ne7����k��ڒ^�b���Y��Vs�� �l�$�@��4T�,L�B�#u,�J�-�O�-p1�ݟ�	7�E�f1`�3�)�>z�#���	���rr9�^���w�b����TQ�q��(Z"d�hM�PO3�4M�	����L��YÛ۔�+���� ���׼�7�0�	��S\bVS���Hߋ���52纥7�?��Қ��D�Ĥ��_~D؞<6�0�٫�J
C��������I=t0\�ht�Ӳhot{z2\�w0^�O������>�]j�㐂���-ǹ�:���y4dD�O�[񏽚����p]����H�s�ТH`M���[�b�H�]#�?�z�ΩK�ۻ���M�V�`�{��s���O
�B��r�Rn�@���d�IK�,NC��Db\�D�=��Jf(�ο���C�2]Geͽ(H����	�+��$U��[T�i�ҽ;�_�3���M[t��UEX.jV&��L�X��������T7|���tx�y��R8��%{�ɓ���=c�����k�l��0�A1��� q�u�������
��� ���9��-�ky��dS�sca��AV0oH{q��sz�n{WH���+r��	E���æ�>|�I��%%U����nz���e��J�U�{M�P�����<����v�TN��ϝ^�mן�Jtq�}�<�7���[��1j�n;-�����DS���؂$=w�YϬ����)�\2��R�ذe���bQM�v�]^I���ڍ�\����5��XC
)9�ar�*�M�$X!G%g���3�m��kDb-*��#�����{�'͌�����0��o����{��y�|~�_d�nfT㐑�f����'��t�����Io8�O��:�
Zs�)��ٮ2F�+��-/�K�&f6��kLm��2���؇M��Z�������3]M�V��{��A��Ӧ6[����:�c���S� ߝ�Y0�
�~�;���!�3��#?��w~\���	s��7T���,�c�^��i�_���o��TL�+7�}mc�Ԅ��WlKI����6��gh�� �)r,Ė��$^�����tʴBO������[d;��ƆȌґ�0�5��	��~X���G�|lYarP���;P��l�����*�����W&7W���"s��K�J�6�YL�[�����L�ЉE���s�&k��; ѫ��A�+q��MR�k�Ю����W��;���Lx�����S�[
��\,L$F���@�#�e�@j��� ��aQƛ����7�`k�щ�-��f�{��}$�Ǡ���2�a�������L�YH����̂��V�'�o���>� J����<qe��O�� ����XEu[S����6�y!��E	z�G���� ,���� �%���3� aߕm�o�� |F֥����	�1�) c7�qA�Y��!Ѷ��u*�( D�
R>�
�*o�Ǧ�s�Qs�B��[z��K��C�+���"�<���1�����p �-C�G�xS]�|&���;D:&m���`P�S�%�pˠ���x��w�tc;�0@�`�dL�-��G��X��G��噽���L5]��zM<�[��F���l6��-�6eH#������� �}�]�˫�	"Ʊ� �{�H1~d��g��P2��v��)+�1���S _�;����ߥ<��л)g=Z[�f��b�ݷ�[�f"d&�R�8��7��i5Iv��rG3����O��U����bW�^�3m�e}��\��%<�1���Ub,�:���{ߑ,�`�0w'� �E����l�}�w���r���+P��"�g��C)ڈ0x!g�t�?��b�Du`�ռ�P=@�&vr@;��٘=f�J"�Q�#�Z����J��_Hdf�M��s�]�"9�Y��pwA�Ԏ!�@Π�ON�%�ذyyr�`� �,�7�(���m�mu��x4�0&Xgk�^��\Q�ѭ�2�0�������QCA��o�#w�,i�8���(�Ζ�P�k�����lW���XRm�Vp~�b���"��S���$'��a���m��0��o ���U7/��\�lu	1�['�O�W���R=	]$��X����񽻂0�	;�v-��L��Eߝ�'�d�%^l� �8Tl�I��֦���M�.{Lڌ�tBeG���=����y�d)[���p'��r�{�o;[��|������璷��J�	�Lj�0��6���E�#�ؔ��q>5��_1��L�-��1a�x��s'�/����c1�51��ݶ��a�-E�C��q,hk��@'�� ��
k|����f�5������=��z��L���-� ���ÙGY؊Y����0��&�'k�٠���a�ak2�_�1������S?�K���{ڞ�Y%�����Qc��Ob�f��9𮃙����� ���a�f�����,��dO����0C���.�a�fԻ���@M������j�QD��;���R�q7/Ҽ�mt���⃩�J���p��eb1F��~P�ֆ�5Fj��<��-�
F��E����d�>���9§�F軹� ´_0ц�^��%~õM(,��G7+X<�&��D-��,SC�>���$��~s��f�G��(���"��W�](kF��ր?�#j��5A���g
D,?s^]]��q��8ʯ���Fg9a����&�����^���@zf��Y��;+�w|�e���|��t�)ʸ�8��	��}+�S���5���p���\Dc `8��h��:�^��_n��R�~W��g�-Ng�/!qX���0)0��O��n��U@Jwd��&��*]��9��<e~��H�9ŷ��z�������c@��Ɋ��c0�J �u��}��e����@��J�RFG7h��f��ao�r��V��m���v`bH��U+��"\H����&��g�"�9�5g�XW�o�
���b��N!��8U��`��J4{���"),������.a����C�J�6��A.?
�"Ա�N�}B�̚k>�ɾ����b��~��Z@w�����QS�q#j��0SC@��=�d�xC��\�{���X�l7
Pc�#��O��9!� ���Ӊ;�k=�o��)R��`Lȋ9d/F�r0��ڂ	���1V.7�g!��.��"wh���\���N%$0�))�Oyi�}���Q@1�����������F@	�b'�����b����xS洷�`�u���tP�އ�Y�[J�Ua���! �b����Us���yc,���]a�\��+�]��rX;)�L�d+]#�7�ᵁ��}q�:��,!Ma$�z� o��3�/�����%���>���2|��Wu���E�����x����[!R#�o���n��WZ����z���?턾]��FÅX��`���݌���'�]B����Խ����x���{�bv[\E�����Z����wkk�r��0�Ha5a�3Q����_����������M��:��.Ev�&�pm7�̤1"'4 �Ù~@�!�A��Z��t�q�=�#}�@xN�0�?�A_!4��i�G	��?��4���5M)�20�#����Zv�{�F�P���T���׹�:�x��9�O��W�n�PVG=�5�jϳ�:c�2}Yx�īvK�����ǧ��i<�9e�cF��h� �(�F#R+6��!f�)�����Ua����l&
�n�Ʃ~��yi�>�0se�U,�V��Ǉ���$��v�.I���ˍR��?�)�����F�����/۴7�My�f���^~���TA��qx6�d��9�r�AZ����T�hޱ� s�z_LV�����p-fY�o#��5Y�����sփ���O5�4������	N�h,����o��_�G�Z�FT� 	�yfn�a�*a{~��k]�猭K8�<᪾�Y�q� �/+�(�470�@�
yQƖc��I,y����B@�Ȑ��rb�Q�y���H��gX�[�'�ӊ�t��%���KS�fM���5��y��;	���
a��Q�o����V��(!!���1$�IJ�#ċ-
D���z����@O��s�|�?%d��1^���M��S�K[=�j1�G1o��{�]x�/DR`�QHMBOK;jp�����Hf���+K�����hs��&��v��%��?;F��l��[����y����a]5���
Љ}��sI�ê��{{���0�Nf��å+���?�"��Z�$��ޞ�{rނ{1 ����P��u~>��5<�4����՟�<s���´T�A0n��娯��M��i�$�6ņ�،���H
��y}s ��C���'�樷�"]��hh�Ts7ZY�����m{�tԣ{E�mH盋Q$o����b�=)t*�DZ@![ m+��-�NpSg�I��M��h}�jT�lRu������$�8SDW)���<���^�>�?���fC�X�1i��7��?;�؛�֪=���ϩ���˃�$;�|�ⶫ(b)H�u�ճ�uW@f0,�璘z���F��E:�w,�cFUV�2�/^�D������������\=�������)���A&�$�F��h$ԿS-��33����XǇ� ��p��<?j7>������Kv�D�)�<7;��P2��e[�a�F4����wWƍ���p�
��]x����j��"t�!{������t	����Hj)9w���_<�K��t�6Z�l��Hs�Q@�Fk�-��-LLr��Xu�s�:%���ԆܠL��I���,��${�R�:_-2&���l.D\�b����Z�Fd�aV|,"w��S��\9f�mV�����׮������|P.����^_�Q�z��k#�������;3��)落->P�TT�(��@�g�ݧ6@���܄��A}ɘ�I]�2���/؂+K?��ݩȐ�8�����6,�2�Ÿ��vߥ͑�DツWXu̷��ھg�yƔ'�}����w���B�g���wa��$Gڌ�t�D��$\
���.��C76�7:��/��o������{,���{���lk�m$�;F�ɡ�ݲ
X�P��i2����L�)�*�YQ��OU'��8�}���m >�g�ܨ/n�Hշ�4U+U�@��;�[:�8�\�\��]2�	s�̚1���"(�bvz#6�ckJrJ��;��ͦ<WX�1�nu��~C�Y���b�(>0�N���A::@$x�ej��R��{�q��J��͛I�ǡ�1H��u��2��3�ұ~���?V���+AIT� �n�nlB7��*l�m� s�8k����pir'�έ̡.ð�g�F-�c@��K�0v�Ο~և���0K9^_D#=揅2l$$�v�-����k#s���j v��_�*��#:�xŪp9�6:ۼ�a8��潢c-�c}qk&�c{��{������N�+��ү���[�^��H�6�0a���.��$CG���y
�@TG5�:�·ݮ�����;֒��1�iR��C^v[�����˙��)���Ю�_����� "�y}��`�x7�����M؎U �D.�d�z_#y��y����|�s�[�t-�z(B���^��h�^`S�%*D�^�rl��EǠe�:���E���/j�n2����(
�f9NK�=L�H�����r^]��Y�D�z�XCy5�*��EWVK��@��<������ֈV� �֪[�QM�Hn�/�Z"'�=L�3��b �����3��:�WC���?���lK:m��~��oC��7��V���.�����X��zb?�>�%<�(��g7�i]y��3���d��>*�	~����i��j`�k��p	MxlVMT������'��pdY��Em��ci9C����/p����ؔ��Kxw�2}p鸨9pR�����}&��"qP� -[)U`ݣ���[���c^7�H"KW��"��~$�Nqta���9�gU�1^�Ց��XlU4�k�Qē���4��0^�x����n�P�� ���yEB������Y�\ WFXڽ��U2���;I�wi+	�� ���������3wr��`w�2%@P�?UPX=��l$�\�ƍ�!����ٯC<�f�?6mc�t��H|h�@(|��t�9�כ�N�@�}�Ĩ:��*̕��c�!���GN\�x�# �Z.���}턎Ň�|�V�M�jl���.�9�&8u�'*���Lp�ɾ$X�q^�m
^`�:�b���èi�3&L+��c'���a�[#C�X��hRpo��CK�vl3�9�&p\఍�5<�;/.��{ ��m'zW�l���%J����;f����G�sZ�&��4Ҏb��uM�+ҧ)�@�x�*�%������C�v`r%O���� QY�J����[B*)w��ph�qՂъR6���1�<u�B_'ӓ�:Jb?j��(G�p��um2 ($gUa�3�	�=;���x%N�����w��Fښb�����Pڰ�%	��Q�i瘑�kdmw�S�lȀe�Ml���CF���O���)R����9�c(j��I)�@��%L8����꽟��P��/��)ǗNPNb�A"9�C���H�0��h��w#����������fp��2�9����bǲ�"h�ދ�����;����E�?ne�mF��G�����8��`5T������E��f��RF��e�ӟ*���[���.N:��p,I�S�����Oy�Ao�*�8����R���Л���gY�a�K�$`BJ�&�7���;� �3�L�Џ-�ͳ(R�IC�o&�E�w_TS�����'>z�N����K�J���ֈY�Զ���|,�y�d3����:7�ê*:�����S�m�ݚ6t����W��xu�E��RU��P-��Uq�����ER�¹Ֆ�du]�\�YZ���ŷ�|}���K�@�}��ō�ބL��5F�����T����,�,����7���19���-��-�/ý?��T<rX8�xB��	������r����p1�(��'j���w��X�:�#��`f;���ߟ�	d[��
��L�W<�dM,<KK����X�qǪ	�IbMt�BL,=��U�2}qjl3(A{�.��-`������оuK;�;���V��{^%�Cd��IJb��*#+�	���Tf�V�%g��F���i�5i�j���_���T'�!�9u����.ID6�r���ʮ%���!�B����&y]R�\"d�=�&�h�m�L��[>�J^�S5�-2�%�X�{D���*��dR���,�SVE�����~X2`�=*V
�����E�OgN�U�I\�R����=�����&ڭ��X��\��������w6�`�bໍ��+W�_���z�ʰY�?��1bx�S��Z���-kU�2��\ܙ=N�c��jt+�{�o��:S&�E�%��7C^ͻ��v#M�Ul�O6��~˰��K?#o���,ӂn[����Z(�����3�R[��X��SP;x�Os�k��^)�Yi��-�Gv!g�icc|��i��ԋ��j�d�O�T%Q�iR��1��-�u/��T:*0�R�M�^y)i ��p
l�	K�J6���di84���yq�z��$W1�W4�t��ip���Y)��tI�1Y������..g��1�ؿ�u�Y����O��a���o
xwş!�k0)]Of3g��Ք/����N�+��$�ɋ�p��dh��X	�)�q��2T���+�~~8[���� �#�|C,�l#����|��?�2"�w�X�j�1���a��`U���E	j�k{�s�Y�@�&��!��B�3����`41v��ɺG�$/2V��|��ӻ����BT�R��>�W#^�hf�)\�gC	��iU���^���)5����4_����,k��/k,~&�:��7<�Rު%B]��VN�6<����?5WE��D�J������8�!�:�m�D�A��y�܋�������\�C�J+�����9��/%�B=�3c�5M� �N�C�:W�C��\c?�=��Q]�W�B���.����.��@��%������gO����J��#5�B��������a?f��*;�p.欨L����1�` \,����!6��Eߞ[�!�C �<�
S�u��b�mkZ�mV��`�f�P�~�ݣ<]˰(��n���y5��,�8	�Ӆ��a�r4�/��+F[,@�).Zp1Kl�dV 
��c�T�$m<j��<�����
��xy�|�.WR��|�we0M�ή����D����*�\���].�+B��ep\y��`6�ٚ!�/�pH?o۪}w�Vu��\��D�<�y2�{m�Ȩ4O���"�HP˚=���V����$|�ΥN!�r#$iw1�7�7K������S(@�}Fa
w���*1%% 2S���(���clŅ���*�
#�;��<�m6�a�`�֤&�J^�i��&�	X�5�t0%�ɷ���~����7�wf�~�LVH�ƌ]Xpi����y����>mπ"}���*Lk��z�%r����<�jl����\Q�w�2�A�WR1�D*R���U� �2�o[��]���Kο$��Z6�?����@�P6e�,jm�éo.�fD����e��]�R�v�(+d]�ދ:�T�� �̰�@K���+r�H�PK����+�������q�P ��<.h
�+%��4��6�"$o�o�ļ!���Dխ^q�Gv�1����溤�Ij6�|��!��P��9��`�)M��o�� q�^_�;�'|�T�ф�"*����3 ��%����(���@d�*�18��*�ǶQI媹���,:7^�۳�𛜆g˵����c�Ƚ#l������C5?O��&�u��ˈ���M$�0�s� W��Q6#����sj(J������N�8^"��� �؀D��uH9�΂-�i%��1�|�d级Q�]S���4��R�@�%|�Y>�z+�u����l�:Ka0���P�{�ڧ�V�����?#m�ƻ�[)�q�IU��B*�#��P�j�u�M�5@�� DQ��r��`I(�n&��N7`DO�&d#j����d�O%���ޔ�hR�p�ǂ�Z�P~�k����=ؖ4��0���-��[�鎒��+��J�31�����5�O�3#���&E���ә��v��&���+�k�.��ՠ^/���롈[�pR��Vst	!Z�x[U:��k�׶���`{g5���Æ���嶒�\Rdu�ZF�MX��.�2���,Cp%��4c>������KK�r�[P[�,�a�:�O}�e�ߵ��N�.A��8wQ?}���� �'3�����E�1F���nm}m`�
�1�LO��-�"�.�G)*��P�?n��JԪ�P;R�aƙ{O9we#�0g���s=g׋�}���|���A��P0���s᱾5�.q�]���5�J����]�D(�/51��VOpD�>�9�mE�/T_^wZ�G�R�_5��C�6{��&���SxM��z�c
%Ta��#us���d�b��l������@���+�z�%���%g���NeV {nkW����'�(�?5yS���	|�e��	Iɖ�9���3�0Y1a��T��a�gx�l[��:aN&��$��d�g�̠8?-��4k7��]��f!���hF��MLT	�B�7��rr\λ�`�;pA�}����"�(Ӯ�2�r���[��M���R��9jB��t�	9C[�Y�Ovb��\��,�G�_DD.�ق��^��Z$b A�Wv����鉓;?Cn��7P��3�ɥs`��ˢ�� ��X�c@ʻe�z&_c�Yw�M��)pj��w0i7�/��^���#U�>��-��2�+�Ea���\H6�b�޹ͼ�zkrLocI���U�%��`���JiH����0�nj��E�~�e���l� М$�?gl�����&����j�_�T�����EW�;��I�w/��j�;�B��g6r҅����ʽ7~VH�^34��m��  B�!O3:HyJr����;��XĐӔ�~G�r�P��;`?$]���Ԛ�$O,���1�.ʅ��Z�9���Y��^w~�e��Z�kH��$ލ)�N��A��7�*��Y��p��2��GhN�`��ys$'�d�aEXZI��E�Y#�w�n�aA�w X�j��P��.d��i�5
.��D��A3��5l��0���X]�"���k~�OG�+��"�f�T���V��~Y!���^�o)�@�Y��˘���h~
wH�zL�52`? �ZјN�P�����'u� �_ �\�)�6�#⡂�Y���v/j~��{yK��;�"��;Y�4^c#d���^_8�l�����#DRԎ$����2��~��1���PE.�<Q)KG�D�.���&9����:����&�{7�R9]�%�V���z�˖Ӿ���R�YR�1���'�M�C��h	~�Jv1\���/��(�>��u��vXi�';�^7gN͍��)ދh���-���L" P�+Y��7)�̓�@7�?�A͗!�
�6�e7�Q�!hg��I����7�[��P��V����,���8��N�(�
�=N�����(o�f6%���[���%T�m>������kʏ��e4c��ѻ����ɟm�{�>�*�/K�*/�mA١B��'�b��u�)�g� p=}�!e�C������ 6�<�׳a��ߘ�?K��
��c<�;#9ƪlgnݍ�wl_�����A�Y,�J�e�JE����7���d&�yk`㑡!��r����pV�� �����h�w�gI�c]�S��#���������	@�h��fK���x^�I���{(�(�\��M�
=TQ�ޚ�j"
A���Y3��Az�L��������@�4\�%S�~4������0�n��{�E����D(@�|;�gV�w>�:��}c,n��*�~۳w5H��P��pHi�f�y"Gד��(�b���jzP>-/���b:P�������3@��AQ�Ѵ��gG�:t���_n4�W.}jdV8��Y��/u�z��D���[�gw��R�%�*Q�2:�UG������͒�k,�(%�EyXE��px���)�KB�8n�Lpj�DG�����L�dd	��Z�
��Ɯှ`�>��I|�*-�(���grI~��M5$��R��y�D�˫�( *�nT{�����qKs
a@��������ϝV�m��0�rE���f�iz�ߣ̠E�8~�P�J��2�S5���G�g�R�{(��0q��^�'38���������D�)Jp�/�g�p��6���)����}��R���n�.�Z��-���Y0f@����[���#���߯?'z<Ȧ<g�>��O���gH�t��� VeY��t�ɫ|�li�*ֿ~e�b¢��l�;z�!H��n{���Bd�k\�>�o4|t8iۿb�ۿQ�!�|�^pr(�������wB71��lr]�j!�O�]�U��ӠiQ���)4y6�>�r��o�#�Cd�l��!�/��&+ �(���4ǥ�_��A�h�8�� ����k�A�d�W��[��nq�����f8x���U�`}E1�{��č��+�~�@��Wr|D���� ����U穮���V��\Rt�����],�'f��>����x��&y�QG�b�QtS�t�2$�S�3�q��:�˹�
�{x�"����3��T��NԐ���%Eω�"F�B���	��*Vs��9=7�� �����2)Z��F��~��r���-���`Aėб2����~��OX���GU�V����~�DP��TU���0ԧ��7�~��/�f�qT��w?!@�n�����|z���@}c����l�p#=�L[r��j~�d�d���K+�+p8z�l�܀���^ڒ6"x�E;H��R+�!M��^�>F�[*K!����/��֤���,���l��C��ט��>�9�^��{),$Ň|#�C1�������u|�LS�J��	e���}��u,7�G��_ISԽ����bL��A"b�4�s^�Z���@�v9��a��$m�ˊ�%rzW[[k1t`�^ \���̹�&��*����!M
�afzh�r�"kJz� ��iO��W��PN��1�ej�Vb|����o�̞0�%�gS�\a��L0����
W���{���n�_�#�p��{���dV�V�����RT���ߐ���~������+5O-Ѐ���9��E3�S��6M������;m��.P[g�����qng6;8;�*v;{��5�������s��uB��tMi��zy�<Ek|=�^��u2�Yb��D�Z���jA����d�;3��µ�x	a�k��WW��
7J�<��i��UYw�|)3��/�KMd��,!Jw1�&	C3��[��c�]*��������d��OF���TԍC��O#%�tL0H�9h��Ĵ 
��Z��]6꺩�~rL+�G�7����@����
#'܋?]�b���]���˓��\gB��"g�We'�-Xn2���S���_�6������>SnM�&ͪY���Q�C�KY4�ߋ����iv}�D���tp�,�$�;u�k<_�_�SrC�_���
����[�]��Ov� �[rٱ�=�sOt	�*�B3�37�������Git=�n Pٌ~#����rZ׹ipN�=��]�vk��h��	�J7�W�h�+X��Y2F鈺���e�-[S��.���=���K��@"[�����0�m<����.Yi�1���c ��q��c%˴�nn�����I9�I����G5fR�^��4$O;��,�?�!���GsZ]ξkf��m���Vd�N�j*��xN�7_�p+��>�9.q������=r�����G��2b2�g�C'��P
+2���.n�)��I�QhM���f��Ma5Ѡ#����^g�)a )��9_#sO�e<Ԭ�� �Iz���˅m�Cx�Yv��{���s�
������vv�h�;���1���&�P;��'�{.~ɎR�r���s|`�EP�2��̙��+�� ��|�h���a�d:�W�"B[%v�J�aD��Y��3⵳~K��u(�M�CΌ>c
2�JS��L���T��-c����U�\ #&�N��ҏ���8n��@[ʦ��LJ	ȓ۸@g�JS�
N�.��C�~<��Xde�crS��n�*�h�������n
	��V�q���z��~���;	�JT�$�,-7`����02݌��a$�=���Bv����g|? �0��
��1h��F�;�Q�sg�*��?�+{Lo�)�+�)HƊ����е�挞,��3ë���ٹ�2�~7�ş� I낂��ak���~��a���iw���pH�_tShqxT�t�Mo�Y�?R��=GJ��b�5wijz��!��`ue09W|�^^�	��wds:�qƓ�hr�[��p5wg��Hh��²���Ty��@��7���̴n�
���'�WڔG�*�Ta�ArL�H��L�[Ψ;g�T��r���}<(4�"�EJTJ4�������n�F
h,c9��Ğu}��^��v|*q��˟���<�y��-۶��(h��r�VNęίՂ�Z�����*� �(/Ma�l�N��I̞Ѭ�]R�/Ў���Z�h.��:�S������Fʙ��[���\4j�ZU;��-OyNQ�<���$���59`|�c�>nx;�Hk}6;����I76F���	�dujnB�5;�$�;6,ڥeJ�>�E�e��Evц��/�j�"v3KL>MK>q*���w4tߚ�|FK���[��~"�'��m�Q���օ�I��]R��y#N���/���A��^���b�YS�ۗ6���62ڶ7d��e�y؀��ZTof��LI��o}�����|N��Vq�pR�sf���oI��tR�U����ogvX��b�l�� d�Lm�� \�F�2x)J����3g��B�%-��䏯ii���@�8�WU�Tq��eY������tc���T�k?�h�%���Rn��}��	rT�U�D!��Ew���[���mq������0�e_�q�S�`�R�(�3�Lb�	�B �㋴��Km�H��d9�6��>��lNז r����"z�}��N��{��(Ԥݡ��m3w������ n�*	n�~��.p��� u��y�E�1��Y:��VP1��%����#æ��U������h�"�M�j�F�.Y��� �g��d�y����N�	�C�ET�t��c�<����;��Y���ڊ!�w>�����cp���v��L�Ҁb����|0�����7�``�t�)�%	��B�?`D��ni��͞�4�3�zڔ�Ek�0�jP����/����Qv�X��e��X�xG&>'���:cp&��g={�;j]�|R�>��>�}��î7�1�\w_���w�>��b;Z����G2H�uy��~�C�cB�JI����p�	x(�� d=��:f�h�|r�]UjJ��ðj��6P�N�җr� �Ȍ�q���0��>�Q�)X^�K�c��-\_:.�FEw7ۋˬ��פ��ηv�'��`xު��g����_d��_WSI�&'`V|m�Q�5-k��>/
����A���b����x�'�࠸{��t@�ֽF�C�=��Bf*=x(����=^'��Z�<���bV�2�`��$٭"~�Ƙ����m��E��bs�s;������-zڱy��#r6e �7Mކ���(��ƛ�K#?�2Wi���F���\w�jQw�����(=�:�u��]��៑���K>�Dy��Άל�����A�h�ȹ������;�:[���e���z�zD�g�q�*=a�H��(	�Q�̢IPX�]��7�R�����hG "�s��.��R���M�6{��{�\q���Xl�lG�Mx��\�n���˜G��i�4a�0_ԝ�Yض�6�'R��)���>S�uJ�8��-zm�eC��ȐfUA���}I�4(��������bc�y!��M��B�^����������K���8��vVSwVG�<���@+yB�`��I��Ĭ�Z6�պ��^e6���E���m2bNk	sy���J �0�F�A�0J_+�[<���������'�w��4ܷ>W�ڌ{â�F�4+��
���=E�5�)�B�1׸��S2)�O��V�mW*�J��Zf��o%�u��J������2"i��<~L�e����.fݩ�Z)�7 z�h3���hk�;Եo��b��(�
���=S�>��AZ$�?$eB��Y�������7'�j�a"��-{�Bzr��Q��klA�F���IIT:YHԮ~��h���Nm��!�R�!��lL���	�uB/�?GP�q��.<d�&�V݌��t6<����R�o�i��5�hҢ/�
@]/,�!"VHg��KB���o�T왧d�6��Ѳ�E���,h�4�b~b�3w�ƚ"��=���Ze�J����믉�*s�7��"L%��k�]O��>T��˕X=���q���Il����D��3�Jy�|�g5B��9�������!~5�~:�ؓ��%NP] �!b
��0�g�%n�H�m�4(Pcv��U�V���ؼl��ޏ�S\��2��<&���N��Y��C�t��G�����L\F��P$���s̠<�!DV,n��C�>�Ȫo��r��푪N6��(�����6��)>���lN���E����7��/~bѬfu�x�4�́?b��Z\��Ѣ�@�q��͇Qc-ӈ�����4N�Q];�K~��މ��~"��2G��g��G�)�0���_=&&��0����b%lٝN��*��P�8Sq�:v��6;�+��򛂦x�U���yik�!������'_Gl��� 7 Ą�y&���:�6��d�s��o�g�xZ���+S�8�%��=�?�P�oK��/�����7?ӎ�jc��/�;��! ��4*��|��{�6�+�H����Y����2��x䮘p=�����(����d�<Շ�)���1��K����a�ή��&^o@)��8�G��>d�����D��z���+���ۂ{K����:.+Og�4{#T9g[ϼ�a��Ñ/�;$;���=���nL���=�GsuRU���g�r�)V�� h4vQ������J������	��X��H-m��l�&ҙ�wㆱZ�C������I�l(��m��?��4B$��jp1E&h����W%�PE� ����: �%�Ĺ��X��=�H~�	(�W��	(;v#Oz�=p�m���/��L�9�҆[]k��{�K��}��9J-�]�MT{���r��hhD�%��PLp��tU<9n�'�f�`�It���C�ۃ[�)�_��3�=�%��4�ĭ����aE_\�⿁ˆ� {�[�?�nI왁�����N�
`��jeٽ�����m�,h9�
O��]�U��!B�@���7����.	�6�������<'�}z(o��6�����N��3��'�q��/3aN
�I�tp	�� �9G.�[tb����*�K|7T	{�
d?"��q�qXY�	�YB ��xk��L���'^�{1aP@QcQDX��&ͬ{��;�58ĂI�Q��c*+7�ayugs����{��XM��Jj
�O9Jd[���iv��uӯ�j'��5����,�;�K�S�+��s�r�*sYp?(O�V���љL7�3o��C5�|����e�T���-�b#>� �vt�� ���1�M5(����Q[��N�1�@�m-e-�omv#�*�-{&r�z�6�u�0_�?)d}�6b[]}�&V?��׷�'.vm�U�#O�r����;zw�ME"��c��͆V�EAgYy{�����-3Z����c�%�����;�/�Mڝo�r��<@B�k���#���ϏlA�����)j�����hhu�4~/���!e���+{��/�z�#��&�xy��J�,Nߢewh�]�u���	�d��pf{�;��pXo��*�f}FA��;L=�CwkxacM��0)[��>�H��ԂL�߁�����6�E��Mne/5+,*PU���0&aR����,�z7��S�Dae-�%u`R �Pg�L�"N�l�=�h��y���ְD��=��[�Õŧ�x��s�oB6�#�DJ���?"���P�.�� [���
��r/��*����ɜ�ˊ������%��o�r����>�$&�})!�p'�_dt���As����w���		�"{̩�b�Q�?.��~�˧���1=��ݔ����xer���W��<�j�)�0����HB�Ŵ�]�٨<��G�Y��!�δ��6r���q�����|��:��4O��qY�������L��D;��԰y��__V�K�����[z{��U�a>X��Q4�^�؏��KX���\sk���I
~��Q���F�6�0���9C��������9ۢ=F|����&as����[Sa'd���E��:d�R��W��: �rC��Ǧ�>���N�Z������lnC��]��2gD&��׷�{s�A�r�,xP��׶_��!.�%De�@Se��K7�[������k�V8�G1G�����~���VR�@Jn��YI�ؗ��'��;��qLOs�� �����_;Pχ�^��W�J\O�E�Z'J_��劮���cN��a�h�M����wh�w��}%�>�� �x,�8� �{�-Hκ ���c׏����]��a޷f���tK�ѱ�C�������U|��_�i���۴C��*ʛz�}79��c�K`��O�)��>>��G5����w�X�
�8n�ޓ2¼��r�!�z�-�z�Hӻ�������j�~k��vkP(�B�?$��vg���{���q"(���|C�M��ԖV7&�����1�Q%��K�Qޛ�Ux�#�̎ho3��E�(��Eq�hiU_ʻ�g �}��L���o�N&����'�){$:8�]����r�̧M�p0 ���9D��[&��������`�V�-[8����#c<^�b��Zݐ�la�@qKN� ����P8	a�1��ͭ�c[�O�ns�W��W9��i��n�m-i��K���a��y�����dG�)����\Ne����r�����o��:~8�{t��Fr�"�	K�%�����=s�;��v�g�� ��*��-�r(99����y'�.?��X�D(Q?��\&b�q�ѐr��8����{�Xz���y�t�E��J	�l���Z!DSb�jY��l��K#m�9������~'?�8�]珱����H������9W/��f�3��r�Ay6�X�v�I��0�xH^�����}� �Zn3a�9���Hٹu~祡Z��YU����>���q� �-VMLV�pݣ�Vv��>���^^_y�0p��{d��)�Q�U$�Tġ�gUm��O ��Y�8D9����C�[ؿzt��8�{�Pf�y����l�ܻ���թ���~}���O3�oh�>��_��˹�Wc��k����o��R ���q?a���8�(�}q�fj6�Il� "I�+�ޮQ�X5�2L�D�L���F	$��]�Z�q6�>4 �<�~EZ����PU���1I����9���<� Z?�W<�����%�A�7�L�I�-|T`1��4o~l*���U���D�5�hY��s-�~k�Ze����8}�9�E�*p�~�k��*��}pFk1O�}�$]���y��-VD�|8�Uk�X�[Y��'�ȍ�@��_c��k'�p�,�Y�?wIe�in�������d��r����4�/0�4�/�ES�cP���5��g� h���E�c@�,�Spc
R�6Y!%8��{qFŶ�|�`03�S��aL%\�)T5��\a���8�n���g�������3����'���Y��?�ֿ�II_���i��P��z�徑"c+�|��nG'���oB�1�0kT����dGԔ�{�?�	�4�-%���{&�O&O���\�Qvf�4,b���t��v��d����U��C��5�@�֯�jv#���:R�Vr}��L��IY�`>;D1򦝂��@h����g���kL���m�`��9�4�;�,�M5O�x��<�N��T��1A�r��0����ֻBN��C�Q~�h����O֜�R��������fzi��7j�.'�P�����A����sE��z$- �{?����y)^A2
�%�X!�<�f��rro���H���Y7K�d��1<��>Ic��{a�6���w�=��)�j����Ԉ��t��K�=��%��n+
80n��&A!�p�3�`��>�U5"�9/�1=�o��7��؂sJ�塕�H�>����U���I�e$/LHMNFQ�&n&@�!�H�P1ZƲ����F$�_1��&����s���i^@�qm�Κ�W�aҌ���Қ��PdC�AP�wC����͙'�/��&��kk��۞�T懗�y�$��ci1�ɇ�:?$ꎴ��"�����Cݳ���s_>��O�b���6�{Ņ�|t�q­@�L�6����O�mS$����FNl�Hu����6I��[b����;J_��G:,���n�RG�T��38 ��|j��V�j{�bx$Z���Ť'���o������;<c��w ^3Ihe�`G�PGCϼ��u��]k�@�v�_w�v��_yD>�<�f�s7b��~��P�E��1���2�|�.D���I3>���$e9�8L��b���ɤw��|З�M08XR����Җ�@�����T�h�#4�S��x�!�������Iy{��O��mo�}O
�:.�[�5?�يBh!�[�H������}���Q���:��I�nè������'�t1O�׋'54��.��"��<�j������)Zh��E�#��-m�%0�FJ�c]k��rf�)�m,�����Q��@���H��"��҂m��Ȓ�./.Vt��rT��m�{��rA��(%��|��م������`x4&
+l�Vz�J ��S��&�:
� \���y��`�8�._Q��������ن���~%����C|�F�E-��D�������T�C��Y�ʬ�jc���%�5l�V*��B�5}��bc��1�r�ޅBk&����f�i�t�p���̐��q��~3i#[M�86�[i�4��K��m�4�t�Q_CM�z�L�e�k�]��Ԣz��~Bw�6���\e�t ��_E'�� /]�
��h�aq ����)������x�&�#NK��T�����l��<x��e��MN`��8�,��#���ۊc9X�&s��5�P����q���Eܵ���:��u�Y9�(Ϸa�k%�h���l�)� {f^��<�>t2p �uQzIM6w\ٞ���qO�>�䌚WS*��Qh�;J�U��+x�8�4����$�`i�H�.��0(�D"�^?�sVJXT띐������?#�Q�>�Q�o(���h�H��Kf�\w�-�������'��DOީ+=HK�vL2�O�ɜa�rq����
��E5��,��}���Ֆ���n\���Xa�zG��sM>���h(�3�S�!���6��/�ڻ�C
���aw������H�5�1�#�(��X��M�V� �� ٬��}L�g��l��� u[�r��K
@*�Mo�D.r�r]	�S1��ѹ��~t��j��1�D�oL�g�)Ѷ�3Y�w�A#�T�4(
kȼn��|j��F$֭�t�ǣ�K��u�]+R�{���5�֊T?��Fƣ/
a�.�������T��@��AՂݡ�hd�D?{}`�G9�h'�Q�����C��	*�� J���������*G���o��-�C5�rE�.�WFDW�II蠟�4�)G̒�"8��/�Js�։Fm��+9��0U=�A���s�z�ea�s�Kt�z?|���V��~݂e���k�һ�h���d*�ܧ�����%���1V�o�649�]�^�4����M�D'3�+��_]j��ǃ0h��:�5
˿��ů$��s4�c����&����NʏQ�<S2��X��dDn��N���!l��?�A�Z)݁D�E�Ð��J�$��S��-��=�X�Tc�j�NR�����XS�Z�2�j�����yY�~Y*��q�JΨ.,sJ�s~N4�O�o	1'��=ff̬!6�{=2@9[%��
�NҬ_}F�i T�
o4N�P=z��i�On��5u�i��(�9���v����:�4�ѭ����ٌ��rΥM���I�Z�TG�`�		�e�GY�n�Y2(�����#�A�v�Y��,0��t� 1��#��U���Q�{��Ę�q\2m �����\�\oL�ٔ�+Ry»��ײ/�!ϛ��
�VU�Kg7�B��M����q��-o��fg2fF�g�G�Sq?�]���URe?���+��G9A�ҥ,^�N6���_;� �"q��~���lW,�S����!/(5��X��c,u��лZ�ʃgSrX.�q/w+�ڎ+Ei���]L���kp`0�� ;dVC��.���c 9x����q��3r������y�d�>*��(BAfof�M�߯�q���G�`Y������HM{|	�'��C�no�į�9�t����k`PZsw�-�<�Qe�#+��"���4ʑ�w�t.�o���ts�k~q�Ql�e�
��q����^�\!�:���=�.��bӁMޭ�Ȭ��_�lR2b�T4�B0ߝeuf�B �9��X�G�m�"�:���	����0�'|G�4M�$l�^�C7���2ΰP�l[,�I��8����J�%:��bZA�B��3�H�ǤYI`��h`��;�d�,�P�n�|ʽ����7�3�<��T?[�Q�y5����D"r&l�<Ԯ�z�ea$��iN[q�	Ԣu1^��j_Կ5ѫ▃ȹ���y�bhZn���˄v�����Bhdz@��E�D�.B��	r�'��EZХ@q4�ߒq��q�j��&<<�/(T~��շvF����SR��?���'
}���V�Ig ��!$�Ao�n��j����@`.���t��߆�J�A2:�~�6*̀�/19� �4aP�X��A����=���z��!"O��u��iT_����/�&��O�$�@�n��V����� �M�W�
h!�	di�U��	��_��m��F����Y%�B�j��W��f�Y�Lݾ�{.�r@��s���¤l2�����C��#�l� Q��,�n�h�2��Ɖ�A�n@{B�^�o�)j���Q�����l���EOOL5U����>�������d��S�e�ړ��P�!�ʠE,=?���i�2� �lD�Rl~~��u�0�x3������j�O�'-#5�l ��"A�I�����y�D��M�ݻx%��"�&ѐ��}�5Z�C���:��E�q�ڹ̂��TB:{��tK#��V���%U/-���T�+�����5:/�AU?V���c��K}+>�̎|�jD��5݂�4gcϊC�D(�+�ݷ�tx�}�J��(g���]ll~)V;U\�N_���������V�CNQ�*d�n�G��2�N���=��)w%���oi�F������9�����{��Q�)_2>�����Fn�7��~�'~i��"��S�KI�x���7$�t�T�]��w+}Hiq�y"�W�E��0�.t�$�4�i��)���0�[�Ҭ��E��F�G�s���b��^�,A����5jC��|Fh�e%��{9��VBbs���X�Z��*��<g��%M��(�0,B�YZ�Z�lz��c����r�L!Z�?��
)�j�Q����q��p�Ϭ�u���N��O��?#�&<VP^;��<��ll���|X��ع<�����V���uZ��YJ!�j�*��~�"Ѭ�?<����J�C��I��Ů�3A�
��+���P�X�2�OXh�p��<�u� �� tt�(\�~sX����_��Xu�j�_gc��_�71�Śd�]Ɂz�����k#��X8��u$��ok�M+v �y
91��Me�����)  ��%�Q.�/SiHv��*'.+R��]ߪp�	��C���v#����e ��ŵfT-������)u��h�U|}@�i�c:�wƐq�e͘���}��11���_W��f`��z;�C%w�Gg5cDt��r�%�'>&�,v�܉�T��FoQ�������O剣QYz��s*�*yTT�.oZ����#�pӗ�w�Ȣ#D��M�4<\��Mg�^iVl�Ɇ��_5�n�j�O#��E6{����1k}�7���,�LV�4�H�dŔ���M�"+a��}q�3��u���L�H�o�7_}�{c`G3��,"�`5jc��g�?y�j�ҒY���=��;��d����CP���~o�F�kfn�dRvY`P^VL��!�1�����f�Q����7UH!~�'|9E��cϦɜ-�23�G�p7ۄ7�U���4d���D8�qv:q�Qĉ8�4U���M����R��>�2G(��5�:��������"1&a5�% �yy^h��|��m	z5v����&FvC�m�� ��M�9�&Z�����Iuy��L�#�^v���W�j���h�ϟ�R��\�g.�%1�?d���Oю���x���X�7��twآ�~����x.ڷVK'a���v}�>�q%>�02ʣ�%��6^�7��X�`-�&�t�.�f}����n��D6f���h��1�+��� �G���jQ�	/X#?V���Q�����@�ZO�k{�&{�U�跞�}�C��+jֹu��ו�f)P?U�W��4\�Y�p=yWq�7R\�<��i��h�5ޥ��*�/'������9�׎��V�����w,��I�c��\3#cz�ˎҷ�w)���n���(�Ή�S�'�w|�&������G�����*��� vi�#�B�M����c�.FH]ʵ�hR�U,�5���I�SH$O/uc�)	�/B4 ΋T�پQ�g��[G��Sn~Xk�'Q�Ө���0�2������	Ò��ú�-��J�J��<M;ʂ�0�o{!
1�7 � y+�DЁ���iV�Z	�?�K�>�YW���1?�w����d,�v��k)^!�c\�GN��Wyi�=��Z<�.�������h�FYh�����ЎHW@�������a�P�/���R�x��:����?,��*Z�zÂ�e���V����n���޹^���P��Db���ޫM̏��K�*��j�X�����}�4E�k4�td��[J;1k�jK��	�G�"�0W��� -JS��RQcɫ	OK��R�Zf�#=�?�XeƻP�X�9/<���y8bL��X�VE��gߚ�S���v1o!ȋ��lS*j�a--�a�es	�Ŝfr,t�F�M�G��f��cE��b�EQY��o� <��ܚd����W3�ԧ� �*���� �5ԩ�2�����-t�~��m �b5��1)/:E#���V�!V�U���,]�Ac��.�e0������}&ܙKI�/�Q�*4���$����Nx~��M�j�Jc��s
B%@q�હ�5}���rN��Kc��u��y��F�NU<L��-ykG�#��Ao#��H %���z.�����m�J:���V��0�Qލ�m�+�%�p)X�m�	Ǵ.<d�Q��%�C�T�L���3La��'��5�Y /%��TEC�E��Y4����J+�O	á���H��o�&'AM�5L$�4�5~F��}2AD��^�{au�0�q�ZV�_�̛��kN;��[�``ꦈ�m� �x��<4z+�&e���{t0u����x[��"+̸����dP�#Xg��F��p������Rѝ�R�h�L���}7]�>V&�d�F���'��`�X tٵ��?C�&K'�C�w�A��Ţ8���:�Q�+�H�do�hl�=a6��z�xB�� QQ�奆A)����dn��B������wZ���x��B�yz6Lk2p���	�<H�U��_�E���t��5� K� h���1>�
-�ϐ���tgK\�����&�����&u��m�a��ކ��8O��q*`���T�?�!�"�(Y�>� w�R�B�Ia�XD,�~
�A���.ϡ����ެƌF��W����Տ3D��O�l�O���iX�)��R�ة�L!�@\�p-��V~̯?[:����"��WE����s#�/(5˃���si�:�Q��aSO��(02�I�p��R����$�8sw(�L��P#�U ��ٗf�J��@ϲ=vp��u�I�_�?����9Rre�|�:oE���r����K�b���{s�Qǭ>#F&_Q��OH[��c��[�� ESi�,�����M���;���*�ۊ�G΅ �o�Ɗ��<?U���pK1�\��Ts��N;0�X	i+�B��Bf;w74X��C����Q�����F�W���fkщ3���>!~�j�����������CP ���ۗc�l���qw6�4 Q#�䳠��^��~z�# 872I�ÿ�;�Ⱦ�W7��NI�Q(a ͷ#yR��� Hf膅�qY����p9n�y69���(AX�Q���N��n,@���)��~0���U��c��Y����o�TZ��4�oQfɡ���L�i�^^�W���0�K�����,�lZ,�7q�a�'��r���Tq�\�N�s�u�ok�n*d����N����,�R}�ѵ6�̤܈����}Z��=���UC������e�ӧO94'�� <��@�4�5u;�q�+���~���P�>���z�g�3N�in��z�	Ƭ)Ṗ�fK�x���]n��C������f�����%\;����`���x�q���/�I�cEl��Ɉ��T�H�:vr�7���1_H�ڔ>i�U�/��),?lO+��7���_Y��<w�n��}��v�~�����ˡb\ܑ����PgWV�A�k����hf�� �6V�:=�/�H�G����q�7�I~0Nk��R2@�=����t=�b��l�b�u���H�I��uk�S��o: W'@��8�(��!8m�tz�x Gv)E�FЌl+��=�����Q���	�"����Я�T�b��0퀾���Re�C�U�fL���lf��g�;Y�R�?yH4̒��?	�J��{���/�My���Q����x.<�0U���,6^�O�[���,�������x��i�/��c=�O<��A/�� �G�fs��S���s�yϫ�_5�^�"�:��ne�xs5�:�/�����;ǟL�/25@�Ӌ�6�*�T�M�D��Ң��
O��&�����n�"l���T"�|��_T��)�:N�T�G�#nແ�up�H�.�R�K�0�O�Fr1~�s��F�����'�������/(k��+H�Ksn��VR 9Kdc��^�CGɟ=�	� ����BE�� �G�~�Gڊ�>��Rϭ�gրڵ��T p2@�:�h:�7.��)!��!�G��о�V�egC�uun�(�OG��ޱ{�0��Tw��c�
�dJEA���;��ƖT��Kx#�xC�J/���.-y�Ӳ�ڑ���r�Fh�����i�����G�_��Zk��R'�G*{^�Q�S@7��F9 ����۲|�)k�6�iZAd�Y�c������2Ѝ��+���]�2Ҳlm<폮 M����U��<B��Io6��hy��@�/�#K���q����@�����Uχ��ИZgY�a14Mp�2��5�������1����������=1���r�`i+	�J�΍�TG[R�[�!�b��r$B�)Y��ߖ��e���oq{�8�E�Օ4�ZSo�F��H�f����2}^�h6�?�J� � \�8����d *����W��#֫2�Ȼf�_X�Aa�{�"\��&g���6`����J�����t[G��X���=P<q�E���T��Y�`,�� �=hZ2�'C��b ����R�V����v(@�wV�q��������[�{o��+�5����s|�j��o�S�F9���y��Δ�t����͔��2u��z�<���i�T�����y̟��˹�C����H=� 0!w�S�����*�Q1ӽ%1�̤Pj�|ʊ����5ݸtEt_��b� KT��Ӏ`�}�z���r�S�ZP�yY	��>�;Y}�ˏV�j���׉֗`|h7gM9�[��o�\(h~S�f�1��=�1mFڦ���NW��Y<w�xz#���K-r�?,��m)��F/�Lx��KE��y��Ǹv{|Z�nB��W�%�Z��4z�.\V���>�3�Kt�� �-o����U��"�h���ūJvV�^��*���܄��k�$ESe1o���W#�D:�z(���7	�d⛢xIO�N9n���o#�D0;ޞ�M��� ��9�|��f/�vBk����~�P�XGOާ����t����dũ��I[heep��� �;H�$}^�>�p��J�aWtr��H?�ڨ��*��5)�4���Š�	�"N5��� VE�G�R-O3�^i�g�H5�0`7Q��)y_����zL��������~hq����e�4����\T&�Y�O�q`ǀ��%�ǽq�h���O����vdM��O�'ے���S�z��&WKq/�G�fP�@�s�Y��jc�ӆ���`X�&�Ǿ��H�(�W#T�gݜy$�CM.K�� ����32��XH�y�ݼ4������1C�F{;����=:�`���y?u�c�&P�����VkO��O�Rr��������$(0��8}ʣ]u� �S9/tn���L�,��?�Fȹ�w���� A��͙,�Q���pG��:{�0��IԦFk�|GӉ�8oY}�6��E%��
���$v��9-:��K��p����m��zP6�lK�`2&���*�2f�A��B�*� s�V�"�0�$�M>@H�J)v��b��oH�;�
�%i��M:��]c9ՠ�5-f�yU��e
��v�j�����.;lk��zb�`F�?�iA3RK��$ P�,��G�5�f/��B�(�B�ڿH��b��a�W #Һ 5���]3uVlfT���>7z�!�kݺ���@��6����m�/-�����=����.���E@x�������_��Շ�ͬ��(������A���S�R����~�6=Ŭ��Up�^!��R<���D����R1;����y$8��X�������%Q�`#����[�1] s�c)��p�1�1
��g��=�j�t�[�����.47��<�	V��0�n� ~�ui�|b�.�]��ب�,K���T�����2
qt"
��r�����A��%k�P�z3�R�%d���VT�r�(�	qOuHP�fN�^̵n��\������!�F~JRESM��"�ґ���[1rΣ�w˦,O��=9�@,n�2M���RB���� }{�q:�`�I:!EU�pz(���t�q0����hK��=}�j�K�3'��.��[��W'=�z�oX٩�\��v�vB���"���B�����w���d���C��sXY3DX��m��)66���� �{����B�~A�v����W��')��i�#�D7� �RhB]��X���ffY�sT���	��A��2Qq1�ނ&'���V^� Gg���J��h݋(��ȗ"7$pLӰ�>ֱǓۓ6�k����#�x*�}U�%�����*��罽&� 1Ү]�"��=O��)�"-����bi��g���Q�5.���E�X�X���<bl]������}7zyU��9g��]CLӒ]A)��x�C���U����ǚ�M>B��{6Ae���*���س@�[+�-�]����ǳ�z���	j=h�e�q�7:]*�����W?�����%�)�v�Q1�~�#\
f�-��چvn��e�Qc� *F�B^�^iv�BYf\�䕦RAߔ�P�n:X�^EӮqN��A�`��*�s4���UZ���y��ETf������(zi�[ސW�Dʄ��u�0��ڨG�LQO��ȸ�c
	�#��}�B��A��{\x���d�;S�9�=r՞����:%��r�I
R����a���؎��.����������~�k7�	�dI��E��܃r���w� �������aJ��1� cRp������F̝Jm�0	[��\�e}�_�r�0�`x�9���^��c�4H8급C�9h0����)ˌ%UA*�$�����}�+N©m&��D��! Y�:+֚�`��1����:R����p�C-A��TtW���w�6��3m��%�wG�~����Y��=&_���f���p�`ݫ�=g��~��0�ms]a�����!W�龜����F1����7���Xk�%��#��'�p� -�m�	�@�b,U�c��."w3���?Y��V1�ޫ����YwRIF��� Ȑ�׮ƒ��8��m���T:x�b�[�|�V�΍w@��AIV�h��AT:�!��Зϓ�>%�Q����#c7)G|އ-#�{��R-v�jU�eV����$Q=*�%��O\ܑ1_x�	tO	�d��կǣ|���X�m�f厐j��r��(���U-8�w ��Vv!+�s�=.�""M�|���b|ھ�LE��t x3(�Qj��7rj���C��Ѳ"J�x��H�������{X�m@����s�?��GmqbQǢ���GÍ�Ƀ$�֍�bt�űe�ٻ�{����g*y9��w�P�m`��Xw���"`�߮�x_9��z.��Y�"�_�v��|ؙ�MW�Y�����/� �Яp�߷�⒯�9/���ϭhjn��2c�#���mf�cjMj�\���p�K�	ئcH�Y��n��|��L6p��ܺ�-��.{؋����ПġWB(�Ƚ~LQ�@�3��x.�ni��q����Q
�E��2i3h���2�I�,?b��u���%�V��v*s���+�"����4�.�Վ�F�E
����V�g�~Z�wK���h�*c����ו
���{d��]���^`��}��*��ؔfP][u�����~=���
*ixT�Z�f��YwYT���^S(+3��j�TǎM��r T�Y�?�7_�n��M��jc6[�*&ҳ��s���	5���3��[�a�ZT>,�����FO�\)ڢ�8<LL�G~J����~t*�f۫m[U�v@'hЀ��:�q�Gg@��A&C�`�I�]�`��0��Xtv`��2�?�Q��@%�IE��g�A��2��Eգ�� ���|B4]Q�Ǹ���e��5z��Jl��T��Pj��P�+�~��Ȓk}o���u���셆nH��vs�jС2��6o�-)bL�y��^�D\��7��l/�+���]Ei�iRv?�&��-Mf�-o\��c��U�ä�(���.Q茀��b d�")W�.�r��i�B	S��Ff���}�~S��q��v�E�%�J�t�O�˝�]I}��⮐
|닩�!)5���ڋ�Ha2#���{5$V�7J:Gm9���1��Hoz�>xrs�BE���ը���Zb�/s�9%��$/�b拉�j���F��IxS�?�33�V��^#�����\m������r�H���5}�Ǒ�(�䞵��w�$��w���bGѫ6�H{Fn�nXB����U �i	x*��o������Ьq�&5��v� �^D���@�A��n\���$��Jޓ(�ݟ\EQ������r��e�i����.�߾:?eQtK����{h0 {t��c����OvGoz�Y>7��m�2������/*G$=7#�|
�P���D�.v�+�(h�e ����p��ۜ�����_��E�.e����6D�gN�e�۟�0f+O�oa�5l[+�k6�#���!��a��dǗ�n� ���!�I'M�D
���`���I`�5p^5��,��X��.Ӵe)��Q%�� {0��%��R*ؗ̄�.�T��O%¿e;��D��e䌎G$�4����'�N���7�� Q��k�����a;��Z�}�0T�0�S�^о����R_0\�L�@y�x�E���)�=���$/�M�i�|C��6R���,�[z��&G��� 8��IcK�����a�#�f	�-���-�:ѽ9�P^��Hh�����L�&��{�7��p6w�+�9��g/���.lkG�����7�׫�rD/u��09p��"XN��q���@�?۳H'H9���n�;a��u,�קQ-�[Ŏ��J�����K?ƪ������7�.�|	����i#���'�����}PBm$sO+U�=�Y�b�VF���V�H��{i�3��\0�
N�Bo�1*YJ�b�V*�p��jG�A�n�oV@F��u���3�zB����~ [E���Gz$�^��y�`8��궍B��'�j�J�3C�+�m��l��G���\@��mM�;�;2��K�P��mn�imIo�E;��]�L,R�+�'SI�SQ�fo�_S0ݺBP���A5�;�(Y><\�s��\�����$s_M9$!L�'<�̗uTA�ےQ�����³���X�]b�]e�%����/o�ϫ0ւO��9�L2��*w�z�r��!�|z).|��/�hDfU������(���A$e���	��5��ο'A�o�^�O|�kE}A�7��>����������Q��ޞR�Wx�\�Xp��fg�؜�OLe�/fHb���d4+��*���w��!�Ho�}Ƿi[}b��~R~%5p�%iΫJ����^aณ	�?�1�8%�*�ߙ˵��bϾ��r� �)�&��z��T�X� Vo�+�1�V�� �Q��@5�����C3�Ց#b��o�M}���(��@�����w���>��>��������\N�4��5T��R��g�"׮ҫD����}������	��I�C ќyٹ_:"\��ʊ&�vᆇI�d΄l���[��u��R�'{N���sT	-[��?k��{�X��(��R~�8_R����_K�j������I�y쎍q�d@��=��a�0k���	͞6#K`K���fCN͛&��5ŋ�
Y��[o�G�%r���������D�:X�R��n��V��v�~��׉ۖ����uO�ULfY��:�"nk�|���*V����&��9mhr��c��&��#�MrZ}��Q�J�RYv�ߞH�W��SmwQa��#�R��$mRl��E͉|���U�rӤ�;�A	���u�s�U6%�\_:��*e�|�*I��I��h����J�35Ɖ3�j�3ִ���Q�og�u�����E�&��0Vޕ2<��(r�4�5�MŚ@�o �%$2��?J���a��KF�b{"X?d�I��Is��a�z�c���p^8�w]+q�O��t�_	f�n�M\S���V����r.���êR(I�$<���Gj$�����Y�!����
�i�����s�%OѾ�L�V�v3z��������޷�uɢ���=�>{���{���r�ۥ�1+V쟙�2˵t&K��.ϼoBǎ���McE+�=^�7|
/;zL.qFN���
W��[��E� �=m��K��
^^��$]�[��a��f fw�#����yl�ߦ߲!=���p+�џ����FFc��%:��=�1q�ؐ��O}�n�Oi ���r6FC����O��4[�8��(��}F���3X�rrZq:0辟B�ߌ��7y�h��"g�P��wCW�դ����,�����:��|nH�r1p�2��[�|P"�K=�Z�dF��yCg��"Q���Oe'�r�M��*`���::�I�N)O����t�,�ս1�]@�v��Ō�l�М��Q4����>M�֍�I�����:c`*y2��٬��'�*	<������r_p��`����k�*1C&��D�"�4�=�����f�ޓ���)�J�2�P��`����9Jg�]�7��+�Ըo�jfM-:ç*�OU�i�m)%�)#�C�n7�ƛC��`!/��*勝�t��bE1$U�\?[����Յ��ܰ Vq�JP�P
�$f`�e�� Ýn�
�[U:�M)��+*���cW F�z~t!E%��hnhxd����Ւ�x� �<ai7��t�<�}����޸x<7|fs�TA�`��<��@����٨泍�-WZ�a�T#����������݉!%�^�k�(ݟ2�'U�Jj'7��!(�<��}�2���ȩ�
�Ӌ|,��2&~��O�a��Z�忄�ޯK�>��/y�f�J���ƃ�h�k@��,�Ǯ����Ҵ,�8e*6NP�b-�0�������i�.���H�~JE+���,�[���T��; �J�$���cO�y/��m�3��*�7Bi��/K�ja��5�gH������*p�@�%�+���P�x@t�~������E��ou��+�x�-X�&�cw�|g�Xr��oe�<��D^�d"�uC����sN�w�ɓrޑ��/0�}�\U��%�	�,�X�?���Bsos*D���uĜ�ޗ[]�%x���p���uy��5���i^��ʝf>:7_ɦ����zc�ńEf�%��o�:��5Ck.��
�h(��)D��;?��6��q��o�}'@���l�VSu��A��_�3Js�y\���(�nS�}4������,F��;я��S.�
vn�����Rց�-�u�	kW��D��ہ�̖ST���Ҥ��Й6s�iU�F�a�eϱ��۔�@XB�o��K�G�d0�CI5�ץ\�O��~�$4u�m"垈ݱ���-�&����ҍ����P5�H��d�ΐ��i>!��9�`M�1Oo�l�h!�������	 7�?%�ڭ���B�Y��7����mŧ|����׀�E�� :��֑�L��N�b���%�@4C8�=Z�� ���S��pk������)����t��emb7$��=JC&u�7��c}�@�E���pv;f/Qǥ�ʧ�m ���o�7�b�E`�td�K���Ŗ��M����􉗧��ʳFm=�S+ߍ�-��ZIq�1G�ܭ���S��>S�{�G�Ju>��z�Ce=u����y*����Ra1�i*���|�`�&�\������E��i�g�e�q��;��ٹK5L*�0"������
~�^kƆ�����Ļ����J��ѣ�_ʞ%q�V�q�¸�ct7 ��n�i�Д"�ɋ�ߴ̀	ҙ����d(��?����kU"U	eO�󾣃M
}*��49]����PV�s.�jw��aCm�I�����R��S���K;Ɗ�=�-�&8jTr/����cn,��d�]��H��8�e5���=�1Vü'�ݎ
|��v�����vxE;Ub�����
�9٨`���Oj`W-�����0{�һY�2��V��g���M�P�,�h
�J˲R+�����m�o������S����$�����M�="��n�����v%u��õԇ���I=�gFv���?B�Ǆ���+FQ�<�5��&R��߁y���F�A
�n� ��id�9�?�\�OW�D�8Ň�{����i7"2�J)dY�٢z4��������]XX������-���ז�)OBn�.�e��-ug�ZQ�X� ���!(�}��b��Јm�!�@���=��+��r��f��$�'��6�c(iLܲ3���-��*,��8not��5w?�������H�s;�#^��@w@s+v�\15x���>���ɶIq�`պɄao��[�K����Y�;.�?n�����~�*5�� �A�k���x���L�f�Nn�v������Hf m�����?3+�V�-Z�-�(���p-ҧ��;P*'k_T�G�[��V��
��d�E��B��u�؜�h(�u�\֭J��;[�Й�Gb3�5\�A�Q�"|V�.+�0:�')"K�"�)��|{RLa8��&����5"����p�7���7��=H��BkU_�݊�[J�(�D�[M�~�]��G�w�k�嬥�P�	��o_a�P;VDӣFH�a�����_�8w���
II:���YL�%�����lv��H��/)鳟���E;��U*ư`�f���D(�J�)�e�ܓ_����aE�q����.�U 1p��cvi�ʨ�+�;�
�X�>���� V�l5н�|�k;.�.�4��i4��(�A���%�ƕӁ;�#E,a���uHq���rR�
m�B^C��ԏ)N�%.�4�BA�Z3S��:�Q!�bBbb��:7J؄����U���֛:�l�l�k�+���Y��:M�v&5q��#ۻ4�ڀQ9 	(R�P���?�>L���xR��#Ȼ:$ˣ
7;��RfꗨAG�m=^ �g�P�L�Q��D@�g�x�*Rߣy�Բ��6�$T`V1��/q=��1�#�q������t�y��sxg�n�>�<�C��+����̎�W���f��w��#-�#� �ّ��y����{y�/T�#�>���@��sP?����}��(��j	����	?�����&V�:���|���Q�3�7�o�N-���rӊ��ۥ�-��}���%w����$���i�࡯r�ڥ��X���e#�-��n�d��h��e�#��5|�NLi�z�SBQ'�&����F�=q����~��!sJ�,o�'���&4�����B$��^�����~����J\h ��g������<5�m���c�!(^�춨��!�D��f�v�)�O��=��$P�
z?��2}gj�	L�eP;��78���xS���?�>I�g��������e�%�(/��B�^݉y�pQ�g��D�d��4�vEmB�7|����ܞ�])0���E�;���%c���1y84)��	�ź��piyN���{���]�œ�"���	{������f&JE���*ӵ�~Q�����O1�g�.�����_xΑ�����o\g��z�N�
A��xs����7e��d��HnpX�C��L{�?Z�m���$Ta.�tkLp޿�m7�U������!d�ܚc�zM�5}&�,<P�����M�ٖ��3�G��H�� }C����_Z*��*����8���S����K� j*:l����s����%&�!�	D�;XA\s`{������/�;�4�*�8B~d)d��2�*�_%�|˲��բr����v7��d�Q�o��>�b��_��~�ه�m��HZJ�6����#��Qw<j��9Ϙ�樽����7�N�
�{����v����O�,tT����O���DJz��8�%���5��8�Dh�26뫉b[�
h/_�N�*#�ͺ���o�L��K`�?4��U	��2+��
�/}�Nl4F	O�xl�Y�]P��ٖA�`t׃.�����/���@����xn'ċ^��D��BA?�6�\�PP�࿠��F�?Q�s�`�&Xa �7�w�Q'-a/��1���+���Æ�{_���ԅH5�տ���D�]W��'t=4�gg���ð�ņ_i����f.�����p2�����O�`z�mX�*��p��
���,�c�FT%��fC_W��S*L�T��5p�:sO��󉜐�5ܷ2�(g�o⟧���#�=��`��5�®��S锹�-�Q��}��n���̩���A�X�����T�y��9<֬Ј×���7h����A녉���Y�Ow��a��r!xG *S�*U�K��Hr_<�k����L�R�u���O>��~�x�z���Vz��ӻ�&G�okcNo^��|�� �TY��I&~B��ݿ�!O�ҏ���,ضL!�B��l#�s�)��O�m���;�2Y�/�����.�be���bAc޹�|����$�ktUa �jֺZ�, >i}M�G>���|d��e5�ʋC���Y������2L=���&7_4/��N����{��C�KC4�Z�'������}��YY�T�0�9�}��3:9rG���5��XF�𭵉*^�^��(z�B�Qj�Cnw��*7��Y�{�A�u�tM�B4�{�f�\��LJ�qD���2��$c��v����	mf���Q�JS�u8]���/�ښ|�@������q�xD��`a�R�2���V>< ��ǆf�s-Q���_݄ }gY偏���u"*�<x���ܤU���\n��]Hg��%MBu�^�xYH�\|��AC|��.��
��\Ǣ8�8s-���J��F{
Dy6�-;��XqxHvF�m�4pe��	CM ��{�������{�88��d|����m�W�A���t\B�_���y5��jO��0�|w�-JX�@~�>�?�x!��G�ٿ/�*��e4�c����t�GQ8�ܛ�z��!�hO}���ѓ���bX��8l�G5&��-+D2��/u�^�xH5?\I�v���RHG��}>�H7ğ�����d(2hq�~��\In�Y�&��xt��;�A���&.$�T][�W����>E7�UWN]ƄΧ1c��^şf���h�T�)xܽ0�1����q�́��W�"�$l��	�㼅)�=9�ɲ ��a%�D��~������J*�G�M����s2Ѝl=�&�����P:E���� �=�e��O���=�Q�C��X1��֝�~��O �ࣶ"s �a�j��]UJ:pmn��'Q/ǀ�A��8&�z�)�Ȍoׇ��=Q��p�������7�?�WI�r�\�v������]�8�>
�PjF�>��BH&��U���v�\V�s�K#R�6��7�	��_��r����0'��rA�k�n��n�3�C3��Pw��ʑת8��ѳ��%_�a9�"�L�)�M��K���8v?D��fk��||�ۺ�-7��iu���µ-�!�Q�kO�Q�X���8��4˴c�1�uh�W�	�.�ې������3��w$;��X},�iǶ�x���~���9m
7��J�}��3F<���O��������p>���H�U��8�_����)D/���O�Yha�.����i({�G�Âem���
A��'��߲�@�V5)Z_�"�DyH1����"�7I���ͮs��O� c�\������K?A����V�����jPXۦ�<\��1� ��=3>��}��6���� ����P������	U/�پh;�|�RmBpY���
;aa<�T�vn�?׭=�v7Y��c`��b
��ٖ�`�6w���d�S4$cW6�kr�Z�u1�
���G��B'	ͽ�Q߉.�&÷,���>�A��yi̴]���� ��V���5�C3�e!�)Q��`_�儇{��GŽ8����1r�p�t�nHE��㪈�j��|�U<�<t��?d��� ��Of-9����$%O�8��)^�B��x�b�-D��,�WQ���_o^�쇃	�Uw������|��*U�� ��9mĹM�L;���.'_��3��4�Rku���ǰ����TVB!����������� ?�$�j 4*k�n�0�k���#��+�:��s�S��j�{:���)�&l+CM!���-:-gp��Jk/�kPQ���6R���Ypmr�/oMq^�����
i���?���D�z,���{΃y3$"ϒ��BP>�T)�����7�����H�ӦVȓI���7\�`��GgD��ވơ����N�_�#�˞L0X>�����W(�֥�i����������'.�Z����7⏯���!`@z=�3&���I�M�>XA���p�Qx��M	� �K���0�~;��M�Bc�H�\D�$DS�"� m�~ۅ�\;�bC�x�t��z4���P�k����}ʍ�)5{�������H�^&g��0��<��JW�b=�%Y��\���>�x����b;��H������1���w]o�f:=e
o<짷�l%��+����e�[1��E8Ycg����2q�q�؂�^�eO�K����jZ�.:�!�qtsn��R>����E��MR �߁T�oƦ��I�s�feq�`&HEk=��xt�>���ީ�9�ď��&0U�pX0d6����V��4��:~M���^'')h�� 6�����lP�[�D�:�Fu������^�E�O�e���f�/\e��RCMv�J��IE��T�6}��kNI�h��O��RyJ�����1�_*�]dzO�	�K���i%*�[(D^�P=����v��d�J�X^Zm�)u�i}�@�ʽ��\w8!B��)�*~���pWc��ʳ�R�0� ��E#w=�JH䍍�I���$VQOb�;��W���ro�t�ᇉFʄ`�A���F�X�m���V+������ѽ�)�(�b��Tȓu.r�j�R}1@>:z��J9���-~h��7gO�R�8�S|c�V�M!u��w��t��4�z&��d�n����A�����y�����x���:��`KR+�N��p�$ZB���L���͓W����}���]�b�y?&����աt���E�jz�=d5-&l�
�+Y�,=yD�po�iC��>0H�v��ҘJ�p�m��3�W�(/��W/�h�ʮ//�[�|��']=X�5� r�(
�/6d֎nh��@�Q�M,�d�\NR#*F�n�ˏ���u]c�K�����Q'¡aH�٨��+�bz+�$zݖ�G������(f�v���@F3�n�����į9	Q&�E�i�캘�bt���o�'<�oQ:ƪ�x�u�y|���]�㩾�*ɩ�x�Ѡ���C����bӁ�ӈv�����HoX~wr-#c+pr�-ܪ����Y��Ӷ�#Y\��6�b͞���}f�LRr��?H�idHVE*��򍌫*���qJa�+\��U���gD�w&����'��K�.r>�mi9���3�;��������Hܐ�ʤ��M�dA�fXz]��Ɗ��N��rY�I�gW�#������o���z�iW���A���͢�HLz���䃟£��.Oc�����	(�?�#IM�Tncd��k>Na�;���>3_G!�rI��W���X7��X"x���ǩ�̕��_�.�x�a]39��P`���?F]e�r����P��RZV�qJ'��B�Yޠ�I����+pWl|O1O�1ጌ ~d��&������W�&o��\� ��cYatk��/�O�(��^K�u�Q5��C-�W����N���ж�
!'S��2�������9�0��`v�Up�R��_N���2� jiqY�_��z@���D��NO��>���	�x �o������g�Ǯ�2y�J(�a� ��t��{[2%�q:��e��)��,b���Œ���F�����Ǿ(6u�u"'��)>2�N��&%oK�q����A����nn��gj_]�����'��)-�ԯ���L0���f�UP�X�D���:���2�51�^�؊�z*͞/!�6��G>���.(tSUf�����p,���<_gC����!U�.lG���Z*�mb��r����	��!ȧ�B�7קEw�r� _o;�vQ7�e�I��UȲ��-OZL8�;޷��=��e6Ʀ&��*I��.����5W�,81�? 2�+��_�<CjF*n�e��H��t��!�ž/�����]����7�7�l�
��NN?��&MB��\�33t1���s�Jm0^I8�ֹ�|{�t�9*3f�Vi�1*r�i���wg�H6po�����-}�OnM����R|�;���s2ߏ�zz�Muv���� ��K1��cO�?���2p$7�(�V/(�+��2ܥk�崙zp�#���+���Ck],Ğ�6l�ڔ^G+���V��)�.�&��1L�"b:L=7(HH
J�g�J"�֛͘1�ϙ<����Sn�su����"�\)�H���f���;� <|��]�p#���U�-D����j�jW���=b0=��|W|��&KxUt^Ar���f�:Bos[Q�hP�J+�yQ������!�J�>��,��N����Z�ͷt"��i�Z�=/!Z��3:áJC�8�k���5ܸ�NT>���S��� �� ���Mj�JAbG0xȨNP|+)Z�����Ə��9�a��4�	h>�Z��oֹݺi���33���:���\��V_��]
L;�ܶ?ϸ�����ߋ�1�`M;�g��r��O_D�-�4�N@��N�ܼ�b��[���2��Ó;�bE���N_��1N�ٲ�51��`#ֳ>2d�Hq��oY&hh�� �mH���y�J墀=K��8X}�Ⱥ�]O���A�\�`� ��r[����3>���Ȓ�`"�ȦUҖ}4q�@�$3�zU�W�TZ��(@Z����W!D!oo��STl-�����
Կ��]8��!w�!��.lL�	Xj$v��Oh�A��1��A���|<g��\������8���Zӌ�=����)>ZĦ���o͵Q'��\�?��3��K�-9c��I�.>���C�؊9?YX�Z�dY��`��@��$�P���a,E�_�.��m�.��g���	�'s>Mc����N��Z6~�a��#���w����g���F��;�M"�7T3�/c �\]����E�9����wj�cS���6��9�����.�̦OYDG�q�7,c�܋���f�WǸ������c3�Wx�����jEW�|��h=����mI��~@��)�T�G|U<�H0���cƚ��dRSZ�d]�us�"�|d�7=5{�Z�gȐUOuJYs��ji��L��|�����"�̓g�;������7"��_���+ӹ�e�P]rނ+����R�#��U?`)�l� �V���]���$E'�qx�,`���)�=ׄ|D��kO��
��>k
&�?K^Fκ)��^��ViO/�8��������!�V����H��̅R���x@�̃�&��U�b�5���v�亏)�LV9-�E�6 -%�k����sv.SS�8��@�P\�>y#�L���ԍ�_��;��̟�ۭ����.�n��^G즗i}�Y��k~1�CE:�Z����k�Ck�n���hԖ|��H�}��ǟZ�P{?3����,B������P�����G�P��w���X��!k��/K��	;h! Ra�}Y��7��d����-nL�?��q2���?}���C\�%N=3���h\�����X`�Z-�t��(�[N�7��Js���0�r����X�Q�a�4��4^�]�\f��9�#�ψ��؉jCH^U�"�*�̣v�$��F0�A�Ј������_��〘���# ���9h��nA�����/���Һ�/��w�����8�X�S�f"TU#G=��9����9��@�����;L�w3��9�
��V��2� ����?�n4�+~��[4��o��,n{�&�aނ�M�wX��9���i�\t+]P+��*,LO��u�-Y!�B���"�=�lY�.�x&s.����Yݾ���:�~�T���H�&�i�}���P�tĩo@�<�ϴ^�ￛ=���d�7=��}�rC�5uU{j��l�bI�S��ÖK����C\`l�S�z�D.2���~� ��i�����C�@�#�?�L�,�wԌ�r�?��!�KT^o��Di!��η�:m�8�^,T-�T�(��F�,-d6�k�*��j��ЄƏ�|���5fW
 M�T���ٚ�L�47��u�_S5+�r�˗h���e�gRU��!6Q�2��6�^�Ǘ��OS��=�;-=����r��^P|���>=|����I��\���	1�E�)�뢵�=�i]t:��+ja]��ib�3ދ�� �>�/����ڻ2k=��G���Y)����=��$���1��:��7�7���Aۀ���;y(v{7f�0 �EY_yz���
��A��,��{��FB$��r��B��k���c{֗aA"����U��MԼCqA�c�'���U�i.k��BQ�{�U�_ ����9�G�Γ��fu
���,N�c��#G��M}��^�SCKX>��ԕ�� uW��].�{(����J"�:n*E���T	{ �\��e��l~��B�N�C����Ϻ��
o�h5�5��b�(l5������}�2Ģ}s9�.=��.�}{�R��ǀ��������
CI#��k�m�J����l#Wy��	\2+�o� '��|9����6uaA�`	a���J >xf戎�ꦉ
��U��ߔg�z��;��8���? �]쓺���#wA�\�/=E�^-=�"9o� &�<�\VB�Z�	&�J���(˷évY�ELG�7%|P��HY �N~�!�HEIv���G���g��Ɠ������>�Xz��{\�%� F>�s�Nq�� ��+�8S�UD}
~�gb��I�����c-��	R�kB-�lH���4	��4��R(��e�qVs�*�7�P���2����mʸ�
d��<�Gosk��i��<ҍ�D�M��&u2~PJ�kc=#ߧ�~GU��S6�yP-l�����������RܩT6����B��7��f���d������(���j_�.u8L����h7B �[�Q��xzl+��/ed0��8�%��[���Q�3�5.�	�G�M�!����E9��r�U�Y8H��>>�{9�`F�)�#!��4F���~��� �P{o�����V}?�����0�0zUK%t8�[�����ݨw�|�M���{��]Әb�/��ݱ�� �����2ڠ�	��>�W�,,$�}�	�h́,���u��1�{uL�� ���w�I�Be�� �_>�у����"b��b�6$��PN�ؚ��'Z�O�%������{aR���f�� ��4��H��o����7�c�-L�ݘ3+|�� �Ҟ�z3�,
��>�.�q1Q�Gp�g[�D}���;q2��q����1�KH`ƴ�� /=m\�x}����?����n-���Dcn׫�����kx�7�R5�Gny��E�2��,�֪I%dɪ�MW|���洠J"hd���"����yc;s�#d���}�?�&���r�2Y�z���b�!��c����5k띷QQ��w���\�%G��J9ko�I����-t���#�A���w�^��`%��m��1�|ܐ�x��X�x(>ƪ �ԀN
�3m��>�	Ġ<B@n�)��*��WՅx(��&�$t��|�s�R�w�l�8<Z�x����m؉� �����OsD�~�aGJ>�j%\ua��Dp�5�%:��� ���7��㨌݌εt�ɽ����{�PF�!10�Q��t<�{�j`��H�/�	���y�F�@^īu��,�ey�����;>���8(��x�i����~�#�����9����D;��Z�㈴e�T�Ox���(ӄ8a���GZe������� 	5cG����q^�xf�t�ܮJ��T���u���)`�u�&4�UćMd$ʤ%"�9�,��XR]b�&&^�}᪛�-�l=����է�K�;�'~�m��ԕK+0e�����(X�{���4лn7a�6[%�B1�Xzm�G�II[����3�7s�oO<��1���W	C�����������kUݟ@��1��B�t���+���&�����,2Қ~0Kk����&��'�u��+#J똩V�ճW��s�=�qTh�#����=o�ҴO+y�dl�jԎ��8���؈t�>���mBo5�˒O�U9����h��@�"e����y��%A��n���VyC�9����*��ss"�N�U�T)ǒN��:ܭ��_x���yܠ�h��=�-�*�uoPb�(K	�nD9#����
Hw߅9�&'V��_�V��X�Ek6�k������gJ���{t$Q2�v�%ztHJ�(�QpB`��O��b�}�T��*��o��!��C���F˛���RBO��h�qJ��+��.��u�ԏۏ�Ӱh���١K���O�{�i�'#���y�Ҳ�¯���i�N�]��?N �T�F>�Dua��_)\t�Ξ��r̜�m䤩)�����D�q9k�e�~:�T̘ �0�S������W%ɅG�ݺ�Y���6I�G�T��F��bL��k�������`����VU�~'��0�س2�������w�|��������x�_��,��_An�ҋQ]D�����>)��3uX���j�������t)A)�sF�@��wv�j�R�i����A��)���[��Ob��@O��4�Mod΀ O�X��H>Fy�el'�������>�����x�h]����'������*ccl�[�Z�C"i֚p��jM�l�LJ���z%�+K7�̏ʲN[�X�J�e{:o	��9;��ev��uyxu��)d��f�H����H �uIZ�1	W���gtP�j����kSm��=0L�M
ak~+3nq�a�3��?���$�0�a�"�2e��~�)i�fVf����	L���;9���|�Oz#��s^��Z-_�3
�8��X�,Iӊ�B� W��_ hR�'�W�j�G������7�R�)i�o�(
>��|�ۇ�i��ϧ����}C���*���Ơ��(��VU����P��;�}�������n�-��XZ������z@��F�Lڀ�z��}��N�'j�:�1���&����K&-?����E�?x��i��ú4���X�5;��Y��7�se���z�A���&?�=���c���e��fa(�8��h��I�:�1ZO�%$u��&�l� �H"��I��*oc�Fa� ���u�>���d��Q�û^�l�^!�6k��T���1h��TDzp�h���o���xG��v�J۠��4|��DL� �|P1��q��l�'�2�b���� �[����7T���٣L�3��3s��E�Mߑ窪6��V8gu��?u�  p3-?Ɣh���N'������
i�5�o��u�)��τOot��~�W(�*,��> u��2�H^X���R߯_�PN����
�-����|&�{oT���aꊟ��wsN���Ѯ/db0������b�
5#������� ��7 �p���� N������
i�[��O������ȫݕ�kK�&�;�F�D,[���3sm����!n��Ton��L�����,)$%Ե�Θ���	��5q0N�j�s�Η�/���=��p�Ps	�����<G+� ����L��/LL�ߐTFq��X�W(��^0s�/��(�[����&��y�_9������}�u��7��tT�)��`tw;�:�[��_f`����{��Qj.��C�VC+�:���L߳�;�릪_`%�Dб����`+A�����1�.g��9:in��J ��Gj�7���ݢ����tvmh�ŕ��ȅ���Jf5~+(!Y"o������Ȕ�S{F�<�Wf�ƨ䚐ҕ'0��U�ç&���U�NՃ;��y2e=;w_+�oōJ�LFfd��(�[W�Ҋ����N�X���4�ǝKu�;F�� ��6�������5n/G]H8[ܢ��ك��j�`��_�L&˄���y�7)��@E8��n��v��"|M������y`[��
�	g��<���0�*�hu��p4�X���W9�|/5C������$HHX� ��L�����p5]%��`N�;��q>I�{�S��:�Y��l}�d�K4*��t�����Y}Q�T���g2u�ί�zQM�Ը� ��1<�Q�k��ڐ��}z�ms�aaJ���m8x�š�������4Y�%�n"G�&���������v�}L>�!"�ח�+�"g|\u��<��`/7��!.4���^b���M��U�RZ���9�9�O�˛#V�S�	�����_arֆ�Qk=bq�S����Gc�6y��k�:((��!_7	R��
*���8��+���F?�?[�G����9��+��'����+o�P�t�r�sEgu�!z6�u��?u0x���Ɇllw�[�ɕw�W���je���pY���v� ��fo@���Ӫy�~}-7�����-eH��=�}>���R٨��+�{#�"�S�"R��jI� �ʀx����b�x�y������,��qԔeIGT(�9wB���˟H6pA��
��_E�f�H��Y�ᝯ�'�ͨ�_U����p��Q�t$��ςy�0�P,��j��~ŢF��Q�l�Y}$r�7���J5��q)�]�d��|ϵ�~<e/*f+�����`*���jP��H\���إ~=;�����>P�n�r�/���S��S�
o�M�'	�自�	^U}�<��N�8T��-�:d�N��a ��
��/�1s���%��ܓ�7FGkd2�*}uc��ցОK5�V"�v���j9&�����9贄�QG]�>vΰy�r�i�F��	n�kY� AjۏFf��,����R�3��i&�չ��7r�}Ϻˡ�,�J�������� ��S��w���_|�9n~0�kn��1��kUJ~	s��i��`cmQs��<!�(��-�P��V3�mCN�j�5#�U�O`뚡r�g�
us�����C�����R�f]m֪�|�O���(.)s`c���ɛ�7�@F�t��Nɞ���l8͒�M 
���Ui� 0��DA�X�w@�ad��SZ�ۺQ	~nB�n���c������{Z�B����!��a�Y��4�}L1Re��j����8=��+�5�[b��|Z�Qr����~0q+a���2�b�^���a/w�g��rNy��q��tg$�'���p
���4�|�@��b �b�����^KB�YV�1ה��!s�1��+dS��t����Yt�f�=<��z2������Is���DZ-=����{"���VZo 5(=n����d�-�b��ΪWQik�#��$��7i]3:m����'F+�JC�/ӯ!�h���?��eʨ��T�+��@�����pP��јV����/����d>��j�;���}�zK��85�,�k�l)�~�����?�IVy�����	 Y����^��W��2�z� ���Gc��l�t����&�����n�b}o�e>+D�y�x�i��R�/�e'����@
�(��I�E���'O.��gd��>�vJ�|&�Rc���@W�|[sH��e�-�j��V&Ċ��+,4������4f����?'���><�Xl��߯c��K��	�����ZQ�-����0�r$"ɥ��z�������d��l�9��U�n���$��5 �b�9OXV�k�[�w�,�Ƌ�?�䏒���롽+W�:�*yi���=�����c�d�t
�+��i�t�����0F��!��&YQZ:0�P�����X���� i �÷���u�Hf����5ܣlr�"��n{�]gy(��l�Q��+e���Z[S���s ������tUê?ue�$��IJ`�6K�dR��k��+,ri�Պ��E�'��"�u|���N����� �j�-*{Uϣս��EkRQ��;1&���}���)Y�3��}i	mz��aN�إq���-�J�?���g��Q��I<�wiI̲�jQ�ؚ�^�\��~����>��%"��B=��o�H�7e1�(����	�4� >B����L�g��^��9���aEwfr�޺a�¯�!z��Y]�JnR���)��g�BҐ��`����巵^[��]oʪve#?�(�\]�=&�v�զ��azX.�p1�ז����!�	��'�;eD�Q˷߂�Z��ܽ 4o���?ǒ7����N��	��>��z�
)і�!.��8��`�����Ϗ&n���?a�<��� ��٫ԑԂ�n&E����,�A����6c�g��f����M���m��&&M���=�& ��^����#��.����l�XK:��O;~�z6�3��� �w!F���;ߍ`������,*c��H�R��s =m�P4䢛�(:C�2��5I �`"C�%}�TL��`Bo�� ���"�MD�ec�Z���;U�>uK�&^��ˌ��Y�]4 ����?:Z�����(sN��@�;U�տ�N�U�m��_���x1t���uù�J�Æ0����$c��Ai}��h�������3�3�G������J�����w)�-
hS� ���<�X�q�q�#�^�[e�����/O��)��f^�X�k_�Qy���0��S�;�V�.�U��ZW��S��?�Y��6����U_)g�j_�xo�>U��_�-��4��Ԅ
��z�A\�L�����c���i􃢍�2u�)n����^+�t�1n���������[�_�A�����"F"y����E����Q]{#���y<�QO��k(��@�_��J���sBtaf�����Ņj�{?[A�
]����mi▞��Pr�� ^zp�JA�-&;?%���ӎ4a� 2ڶ0����#t������"{s����G�/q��ϧ!0��8K"(_<~*��8��.��AS�4��Gk"J���t�X[�������S�
.*Xq�Ӛ4��O�;u ߯M�G�hww'hC��K�Vi�|�I� k�W�ݳ�^b�g�1J�c�D�w�A���#xq��2�{I!�$��|{'Vָ~�����G]sU/rK�i��!��V�v���e��-���#c�֔�#6F���Q�<o3�P@ر���p7&�M
M�L�.��E{���Jm3>S��~_'cGr��,�f��O�7<=Ȑ}w��Rs�=��?9�xįh\�O��`V��P�;�0�5M�A�ځ���neu�W]���])����}�<�W*���V��"0z!d� �[��|y��G�g�9��~�/B�EEٴ�l�O:�=#	ͻ���m�i�mU�Y��Cq�q�l��H�"޵�Xȩ��>y��Kq�x��֬�}�Е,-,baq,*Rm!�@D�e�j���P��z��	xu��Qz�g���/�F�������^���t��C�
�-�A|j{o��i:
D�I�0�EeL��5x���'Zǿ`����6��L�(��ҁ�2��>i��\�ѧ޲y��rtw��"�"���A�#�M闐"Ҋ/��Xs�T�E\�����1K��Z1���	^p�6� A��z�~<[�(?���(��SA����C����T���zľu�� ��H�q���Fe/�_[�&F�ڃ�����4BP���s��Lio���58��B�.e9�L$��0z�ۛ���ꚫ�gʡ�W�	K��f:z����P�����W���i[
�C1>�Hq�*�%����?H�N�������Eem�4����<�cDe��+�Ɩ�mm	t��k�Of'@�a�m��c[���Y�ؘ�1�ѝ�DV�93� .�:����ZN�y���$�éCQp*^�y ��?�@:Ώ��
��4�vފ<N�UiC^�a<9=��tjVcZ��Bgq,Ou�#ǿl�QI9��H� r҂�'�=�� �C��܈�U|�Jp�-D��z��1�_A�ͻkD�ߊ��GH�Ra��AE���~h�ε�����jg/7�gD聢Mo�����,G�i[a�ՙ����ĭփ8c4ڏ>�m��(����el1�E0@�s���6S�e��1��WMg�u���>��K�o6�����W!ؿG ~~�����k6,�Ԣ�0��u���"��@��� =Tn��<E��9
I�3T�1@\�L����.��O� A�AA�;��G� �vϕ,N+EoN��$pM��Ť��C\�u��Q9nK�����v�p�F�͚�.���a}�Ӿ�̻ϵ&���hH���ޣ��c���[�w��p/m'�6P���-�Ns�̐}�p�0oG�U�p���ք`���zg'&�7�m�o�Y��4�y!�W�E� s�5rVCX�[)Ć�eej�T7����-s^����pa��@ʑ-	�6���)@�#����Y�H�0��tGPd�Pn��F�Q�]K6��{2.Wf� WR�i�jZM��4@�:3q�=G�S�W&Qq���M��~&%T�[��ʑ��_?��������p+@��WE�jE17�K��(oZz��')�Z&�D�6b�D^������{��LRg �0���>��t�U�8�/50�b˻l/G����x��
�G˥�N ��Բ������a ���'��,$�l1�@Ǔ��O��=iqۘ��%{*���M���q� �bD(��^�%�/XW���C
������"-�?Ƌ
�U�=)�*���,f�.:�K ���|$@�\�;����'�P:�5�A�"c(��y�y3%�:�#�Qzq&ۣ�N�i�� �W(��a%�w�ߠ��DUjϮ��nRm��nw���4����L���vܷ_��b�Fs�ӳ���*�0�X|S�NF�@�}�_��f�2�na�!O�Ʒq��>���>1H2�}���i~%u��)D�����fP�)�׬~�8f_my1����/�l�݊�$i��kH�)���%rW�e|�k?E7���t}�!�Y�� �/Y��7фIo	�h��K�M:o�l~<��H"�5��r;�gF��V�C,�&K��w8ҭ����'
l���7�O.�:�Rp9�5��M�Jċ]�^�t�q��/Az����{���s�'M�n<g��E��y������HHL����e�ڙ�o�'";�[�]��cF�d,��G��&��%�������nV:'�}��K�����y�-�Dʬ�A��iM7[��S:P<�,t�yƢ7���1%ߝH�7��~9G^Yg�,�}�����g9^'�Ίsq����B���)D��1�/��$-�*��10p�V���o�hh3�rE\���M{	�~EiS���^Լ6.��2adH]�~x���T1&�S7�R��>�G�E�ck��f���s=ٴ�rn�I�2j?���iu�P���,�L�QڦC��]�����c�	�s����@�Eg��Q���H.�����խ\4_*�e���7�jO�Dۚ���Xs��V�fR�����k���P���m�=�%�Q���S��4�h��qzq9;S�5taN�l'Ϝ%I�o4��;�q�O
���G ��^�X!zg,wJW]��C��~���.x!�|�(Ӣ+3Y�����X�#���R�����Q�2Q@���M�G(۪Hh	�ό�^�6��QWT��R�:1�+���mrU�"F14D"S ��޻��$��Sw�����_3����m�oxh���}�
���7���r
,�i{ �v)U��c��"U�sϽi�a	9�%��@b���9Y7J� A�T��j c��&3�au������� ��ñ5��O!v�Ȝ��%��`�R�i��=ѐ�~F��a i��ePa]m���ya��w'�����"��R��=4y��W��-���Fb[�K�ڷPQ�²7QSU���ύF=�����|��{�5�|���*̃����lTar�ja��/�5���
��S�����C�e}�1��Zޒ|}�%SШ~�5�u��/����6�o����g'�0_��byg��^������Y���LP����nĺ��~�������7��Wz��R&\`{�1��������<��`{��%0?�b�Iϡ�+��=�#�	M����2~��a�|��
��F���UP'Cȓo���s�:Z:�~Ն��#V��u�u�������W�������]�и��E'c�.�)��"_q�e�Px��<�v�	+N$��g]T)�>؆n�"�+�i���?p�@�)��V��gǆ�æc��֗T�qA���	9|���U����2�<�)C����-`��А� )}���QA��4��X=�mN�8 ���x��c�`���x|%�:6=��cxk/M��Q��|�kE|*d��*
�	(�?�uy[���@�P-�w0}���0���RZp�7�y�hs2$��������T�8y�n=G-���Ƈ�i"韹Vu��zZ?�h�o�߂s~d:
�
^��F�>�RCu�R/��c���c��0��U�,8����)�lRm��dOГ�tK Y�|4FG��tS������ያ�};jQ0k�p��.�C�Iy��f}b�w$4�{���|��^��+�Fڋ�}��Б��z�S2����G����Bk�6�&����ǎ��Zҝ��y��-��hǀJE�Q
=�/�u�����[����
^��Y�f�T�	��ǙV%�S�r�;�$[�@��?�_v��e��GG���������M��M^��OC�ˣ�]��Т�jo��\�}��5UHL]�Spu�قS�}"{�l��R���*&M���0��ą�6 ��;�՞DK	Հ����}�+Γ-��6kȡ�m����nhu+c��u�˃G�|(���;�4奏+@�G�>��u��@����K�hSa�����;d�Y��T�dw6���t�k�@��e�ɮ3 �g�4���4�m��%� �����_i9�(%I�g�W���b���Kw礈��D�q��&����*�m�ސj�-��u-�tp.�v)v���[`JF2�g��,�KY������e�OU�>�uoVL�	]���px�](^>Sӿ��!:ƈ.�nWh�.n���9`�X���|�x7�Me| �`�;�x�b��0��!Rr���\�Ө^)�x�����K~)ׯ����Wx>$.	K�*9��T#����I��*X��/r������a}vxwƉ��czX/�/�mݍM�G��m(ԡX��b���X�6��m?ydR�����5�z�Od|"�#ε�(!���6O+E�-��4٥�	�{�^�c�� �$E��,�NTD�M�t
�i��t��K��>97e�9�O����˔�<����N��Nݴey�s��s<8+T: �,[��p�}����������,�Ǳ>
T;�W���<��(	�6Bh�n�L�&*`%���5���Wa��K]1�,\LO��'�9-^9ē���)�%�~���<E&�C䇛�z�P�8{��)�/��Qz/��9�zQ�f�n��h����h{U��=�ZF�Y�%���	�y�(2�a_5v!w����.���)��^��?{�C̏�{ b���ͼ3DW;��ᔷˡ���U�>�_̺2r�0\�k��'ޤ%�%t5�A�7���N8Է��߶"y'�2頙�<I;]Ƹ��f ���#!�<ɷw:q�:�]�g���/L�U��u��6ϟ/(g�at�=�׃����o�/HJ���A����Wy`1�K>�T�h��՜�ň�P:�����ۂ�
�af���װ
�be��un��>\=�ؾ���Y�M�p�������kH�)1�j�G�ځ��C��Q墩4��Z^G��e�^�����2�r[��0t{�ف5`za1�>>���0���n����37�\pk�⻳����ȦS��+���N�F�9bxH7���D��"�9 �OÝ�M%�1�+D%bmb��8g�����y�OF���1L �[s�m�0}B]w��*��Ƶ����+�+������P�@���\�sZ S�IWmB��')�DЩ��1���ӄ���M0~�g�mIf�X��.��z�)$��G��_�Vv�U=�(A��'!�F�}��5'�t@�X���	wwɏ�H�w��%c�����{CZ�4���9�E]L��8��
(J�|�G�׳�<�;J~��EV�C��i�Iq:T�L��h����e��Q@FG���^}�e��*�G�ӑ9�]���l^��X������#
9ڗ'N��`H)-^C�	a�K�LH���CJ�'��Rx�yV�i�������]�Y~*u�1�)�MCD̆��uh��m�u�<�q1���Δ�{*�$���PH}$j�Ot��N�c���vt�3G���enN?�T[l�`�����s�,�t�+]���2١����Mvt�`ۧ`UCA��~���t��yfu�ЖD��x�;a�������;��eJg]s]
�����!Q-��7v�+�6I,���w؎> .��,��k����:0�����������pa���=K7=��BEZ4���>V)��з��9�����P��cҡ�m���"��������@+�� \%Nһ
l����#d�&��]a�0N��|U��o�l2����.~e'q��&�Z���SR�aɸ?���vbS ���F)�����txw]� �����忇��Υ�w_� �>���At���OG$�t�b�CF$��0Kd;��5���@����_P�6}��Z�!�K�E����]�.���JL�����miV��+��@��!N�n{1ݶhZ�;U�fPШ�є�5�*|�9T[�|6/�W1�)g���j���NY!�J���F��������`-��l6�0û��n�ĺ�*���8�8��'� M��"3ʾ H-uD*�]�:�q�7z$lAx{F��-�R�'Ӧ�����hi�K}� �{�Y����,��
�?9������k�9�M�ćw�6Q�!�L9�TJԶ�K���� ;Nd�>�� _��;.��-LZ�Ɓ�0Kh:ƴ��f��E�6W�+w$X���>V1����e\���x�y�5i൯ �͡;������v�q��cm2O��I(�4����gX��K���4�	"�;%�; S�뇈��٠H�j��/+&��hѶ�'x���t���@6�7@���e
1r���e�A�����(���5��0Ž����x�?��e�+Q�Y��<�.࿢�%ZaEU&��͌��I��9.5�@��G��!|Yw@R �����t��=>3G[߄})�'!#��o���v�%`�ɬ.6�@_)�8��enWo�	6�y����R�P�L���@�}�Kk#B%�x�͑wX�7�$�d��T�4���%_�YL_��U�)[BK���D�g�^������\f	��5]黌 u�`��F��;e+�o�X1�O�� 9t9?M������4F��"� KlY���ci�h|�[Sv98l���u"&�3��/��&�����7�z}��e�����TW�1��V���c�����@�m.���t�h����c�����RtO�~�m^�(�h3���pkL]=3�I�Huy����@&�wS����i��	��6Xް/�q��L$���>�0򳑉��P��-���&�r��Z�`Y�*EáN�p����p��d)���Ë]֡�\c:���F�Ư�������Noh)+P���գS����-�
�'&�A�����.:R�-�F����(h���(���&,)�!����>�nر���\
z����h����1Ae�#T���bl�}k���B�����R:1f*�9�z����a�����-/Z��{�����5Ӛ���oc����H��y�{��5���zc �4��lR9bg�AٌJ��e�ޠh<����'�����2y�'P��E��T�vA%��p��j�2�#�P����TA��/}���3���ս�?�s/��#pɴ{��� ��5̍��࣯�VQ��_�[�B�ݝ�,V+�]{��{� X�Y�,#�N��������`X]t<?[�N�
��3���Σ��?@�p�(mx��]7mY;����'��Qt�	{�ߙ��<�&��؋s͊f��y0��t�2��Q�PCS����W�H�>T��q�q]T�pgS���p8�  9⵫ԟ��9Dȥ��-W*h�Q�]�����j��%&�H��$Q<Vؤ�\�p�qO9�|��jȾ��,5�o��аfpE-�;r�a]n�[��3FbĤ��Q�~�q��Sfs79�-���]��������c7J8�y��+��o�[�]s<��!���@���F�#�$0�2O�6�L2���E�Vn>1�H��m�YDi���u������<�����;�Ɂ�N0�.CF�{~�2�
��'��eF����ᭇ��>Y3�(c���\�)q����E�z�;Lc2�-���s�(am��]����:�����w0b��?.���%��u�Jў����Q�zp;�p�(p�¼��&�<U��x���xp��H�d�����'�Ϻ�%�K��|��c�|=���m+�(�UOW�~Fh�e�u,ީd�Fa��ϿDHs<!�F�.�:ˇ�kX����p��
F�_�Е8��-e�����Ό�Y���  ](/Qӏ�6m��J��y�!攷�8��F͏�.� �G�·_���=u8�� Tޫ�q�m��d?��o!����/lu��캼�;�|�D���xMzi�%W���H`C�	�DE�p+ ���� 4yM�lH8��D�Ӕ��b_�ru�,�mB�h�DCd�g�N3N��[�"`3'K�Sx8L����r��zQO�*�C*"4{��JtOw߭�aLS���3)��O���#����r��ę��e���iֵ:YK
�F�'|"�&��؜9��#j����\�lz�F�z#4�a���8��4��.k;>�����r;��0� ��q��� }��z�Dx��'�9�J��Y$b���3 �bȪǵZã��.�m�N�b����8�c\���H[�qU$��}]�'���Y3do)7�0�Z�p���o�� ����JLA���K��g��ڐ�!f��/H�� `Ww�"Iv�YƎEM�:+R��&J63?e�Hu������K������I
n����5���5�4���{�$��b�>�zi�E��vT�m��5r�rdR6�|�n�íE��mFH5+�3 �'��
��-k�8������z��X}���rS-�TstRI^�41�+�����+Eq�ě��cS��#��k��sx�s����YP���� '�˽�HVS���RX����"����88q���V�#j��$��Z�5��=�qZƤ���eKBHcG�!��@H �`���'�X��X��R�"��@�ʛ��WOj`�4<�Q
�תmT�����e�̔�~`�]꒱����{�.����J��bt�����Y�*"��Of�@I �ǬA�bo�*�yfx��N[���5��*(j~�d��Li�{��= ��]�N���$�#.�SG�C�2�mЃٶ<P�������u���1�3�z����.^�O;WDZ�t��Z蔵�_���'�|f�k�zSk�_'=��L�����;s#t;A6?H@=�?����8Z���*f��m<�H����x867	N}��9*�(��' ��579.=, �(瑺%`pm�-���%b-��$�~RK1���J�\��Y"�9m�p2�0��&�U��бI��sW�&4)fc����!\أ	ע��q!��Vt0�ד�A�x)AYN$f3$�4M��U�t���	R��W�{O�r��ܝ�p���KɖCKi�V�j���|׵NS'�H��Q�Ug���G��1��!��< ����ܯ�KNDw\9���5$⽿aSo��"c��o���>��uג�g<Q`MD�8�_J��Z4ؓ?IPh_�KvrŢ}}�>'<�G/���a4���}�v^�O��W#�W͊A���Q�+g5��H�A��_�KuE�C�Z�1p��	�<��Kt�y����m11�.]ϕ�(�D[Q�N+߸Ma�z�{�p�t}�H/u�?_KN�i�Ηd�� ���(�,��Y����:n�^;�MW%4�i�b�ٯ�İ+�w��$9��k��	d o���B���A�̮�bl7\��\W-(2��A���9���g��[�����M�� 3jQ����$�7ApaAи��b4�`�)e�fˌt�Z���)�к�}zgbT�.�u��� ?[�J�۪T�J�� ���v�'��pE�4�9����?��y]�_;��)��e��C�Ҵy5n�t[<mN�oV9�G��n�����bq1GN`$�d�rl��м�: )����Q���%���H��J�Uy�S���3�gӋltlY��e�{�	|۷d]�	8OH�@ui�:�I����ʫ���
�_B;��e��(�uC}NY�����|�}%� cp�Z\Ap~K�����	�e���Ǡ���&�C�	��⧩<���oߔ� ����~���|RVPerJ���K|�l������6c�^V������%�3?=�¡m;}(��q]�._׈���;ٗ��K�)� �D|Js�����m̄�Dp�mO��y�Y �%"�&1AOO}��@O^�r1�HN�y8�ȆIs��c�i�
�sq�R�,����3֝���$�g�jһ�)jI��b����E� 7x����?����덦�N��}�� ~�Jg5��Δ�+X_�K"]d#�z�j��q6�r�Ui���#��8^F#�ݭH���GĶ��a*&\?���]�hJ]��A��5�R���8vF��1}�r�{E��\,�s5�H�F@ƢC�.��M.�Nvx"��Ё�U��P���l�~U�N�T[=Si�X��Ӷ�rn�-�����=l�~�y�|K�w	�'�=��>�a�A�����r�#�<i��p��C��	��5ei"�/�5�w���_�ۃ������#��P1�F�o��,�z�'��p�mb��
�����!p�4���LT�	�s���Ob�����sX�;�|